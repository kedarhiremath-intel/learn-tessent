//------------------------------------------------------------------------------
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2020 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//  Collateral Description:
//  dteg-upm
//
//  Source organization:
//  DTEG Engineering Group (DTEG)
//
//  Support Information:
//  HSD: https://hsdes.intel.com/appstore/article/#/dft_services.bugeco/create
//
//  Revision:
//  DTEG_UPM_2023WW17_FV_1P1_18A
//
//  Module upm_cbb_control_2_cntrs 
//
//------------------------------------------------------------------------------
///====================================================================================================================
///
/// upm_cbb_control_2_cntrs.sv
///
/// Unit Owner        : dft_build.pl
///
/// Original Author   : Auto-generated by dft_build
///
/// Copyright (c) 2012 Intel Corporation
/// Intel Proprietary
///
///====================================================================================================================
`ifndef MODULE_upm_cbb_control_2_cntrs
`define MODULE_upm_cbb_control_2_cntrs
module upm_cbb_control_2_cntrs #(
       parameter THERMAL_ADDR_SIZE = 5,
	   parameter OUTPUT_SIZE = 12
       )
(
        input  logic            fdfx_powergood,
        input  logic            update,
        input  logic            shift,
        input  logic            capture,
        input  logic            tck,
        input  logic            si,
        input  logic            sel,
        input  logic [1:0]      cbb_clk,
        input  logic            clk_debug,
		input  logic 			power_enable_hip,
        input  logic            power_enable_prev,
        input  logic            iso_n,
        input  logic            power_enable_error_prev,
        input  logic [1:0]      clk_in,
        input  logic            so_out,
        output logic            power_enable,
        output logic [((OUTPUT_SIZE)-1):0] upm_address,
        output logic            so,
        output logic            power_enable_next,
        output logic            power_enable_error_next,
        output logic [1:0]      clk_out,
        output logic            shift_out,
        output logic            update_out,
        output logic            tck_out,
        output logic            capture_out,
        output logic            si_out,
        output logic            sel_out
   );
//------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------
//______________________________________________________________________________________________________
//======================================================================================================
//
//                                        - PRE_RTL -
//
//______________________________________________________________________________________________________
//======================================================================================================
//------------------------------------------------------------------------------------------------------
`include "upm_dft_build_macros.vh"
//------------------------------------------------------------------------------------------------------
//______________________________________________________________________________________________________
//======================================================================================================
//
//                                        - CBB CLK -
//
//______________________________________________________________________________________________________
//======================================================================================================
//------------------------------------------------------------------------------------------------------
logic enabled_clk; 
logic [((OUTPUT_SIZE)-1):0] upm_address_pre_mask;  
logic clk_xord_0;
logic clk_xord_1; 
//------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------
//nets definition
//------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------
//module upm_cbb_reg instantiation
upm_thermal_cbb_reg #(
       .THERMAL_ADDR_SIZE(THERMAL_ADDR_SIZE),
	   .OUTPUT_SIZE(OUTPUT_SIZE)
)
upm_thermal_cbb_reg (
        .so_out         (so_out         ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .fdfx_powergood (fdfx_powergood ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .update         (update         ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .shift          (shift          ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .capture        (capture        ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .tck            (tck            ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .si             (si             ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .sel            (sel            ), //upm_cbb_reg::SIB_REG_CBB_REG::input 
        .shift_out      (shift_out      ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .update_out     (update_out     ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .tck_out        (tck_out        ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .capture_out    (capture_out    ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .si_out         (si_out         ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .sel_out        (sel_out        ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .so             (so             ), //upm_cbb_reg::SIB_REG_CBB_REG::output 
        .power_enable   (power_enable   ), //upm_cbb_reg::TAP logic::output - MODULE_PORT::power_enable 
        .upm_address    (upm_address_pre_mask    )  //upm_cbb_reg::UNIT interface::output - MODULE_PORT::upm_address 
);
//------------------------------------------------------------------------------------------------------
//______________________________________________________________________________________________________
//======================================================================================================
//
//                                        - EN MASK -
//
//______________________________________________________________________________________________________
//======================================================================================================
//------------------------------------------------------------------------------------------------------
logic update_ff;
logic en_mask;
logic [((OUTPUT_SIZE)-1):0] en_mask_vec;  
`UPM_ASYNC_RST_MSFF(update_ff, update, tck,~fdfx_powergood)
upm_2nor1_gate update_nor (.o1(en_mask), .a(update), .b(update_ff));
assign en_mask_vec = {OUTPUT_SIZE{en_mask}};
genvar i;
for(i=0;i<OUTPUT_SIZE; i++) begin : UPM_DONT_TOUCH_AND_CELL
        upm_2and1_gate DONT_TOUCH_AND (.o(upm_address[i]), .a(upm_address_pre_mask[i]), .b(en_mask_vec[i]));
end
//------------------------------------------------------------------------------------------------------
//______________________________________________________________________________________________________
//======================================================================================================
//
//                                        - CBB CONTROL -
//
//______________________________________________________________________________________________________
//======================================================================================================
//------------------------------------------------------------------------------------------------------
//if more than one cbb is enabled -> mask clk out
logic power_enable_error;                
assign power_enable_next        = power_enable | power_enable_prev;
assign power_enable_error       = power_enable & power_enable_prev; 
assign power_enable_error_next  = power_enable_error | power_enable_error_prev; 
//assign clk_xord_0 = (clk_in[0] ^ cbb_clk[0]);
//assign clk_xord_1 = (clk_in[1] ^ cbb_clk[1]);

`UPM_CLK_MUX_2TO1(clk_xord_0, cbb_clk[0], clk_in[0],   power_enable_hip)
`UPM_CLK_MUX_2TO1(clk_xord_1, cbb_clk[1], clk_in[1],   power_enable_hip)

`UPM_CLKBF(clk_out[0], clk_xord_0)
`UPM_CLKBF(clk_out[1], clk_xord_1)
//------------------------------------------------------------------------------------------------------
endmodule
`endif
