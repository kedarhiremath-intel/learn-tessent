//--------------------------------------------------------------------------
//
//  Unpublished work. Copyright 2022 Siemens
//
//  This material contains trade secrets or otherwise confidential 
//  information owned by Siemens Industry Software Inc. or its affiliates 
//  (collectively, SISW), or its licensors. Access to and use of this 
//  information is strictly limited as set forth in the Customer's 
//  applicable agreements with SISW.
//
//--------------------------------------------------------------------------
//  File created by: Tessent Shell
//          Version: 2022.4
//       Created on: Sun Oct 29 23:51:19 PDT 2023
//--------------------------------------------------------------------------


module firebird7_in_gate1_tessent_mbist_c1_controller_assembly(LV_TM, MEM_BYPASS_EN, 
                                                               SCAN_SHIFT_EN, MCP_BOUNDING_EN, 
                                                               BIST_ON, BIST_DONE, 
                                                               BIST_GO, MBISTPG_STABLE, 
                                                               clk_clk_bbm, m1_inst_wen, 
                                                               m1_inst_ren, m1_inst_adr, 
                                                               m1_inst_din, m1_inst_async_rst, 
                                                               m1_inst_fastsleep, 
                                                               m1_inst_deepsleep, 
                                                               m1_inst_sbc, m1_inst_shutoff, 
                                                               m1_inst_mce, m1_inst_stbyp, 
                                                               m1_inst_rmce, m1_inst_wmce, 
                                                               m1_inst_wpulse, 
                                                               m1_inst_wa_disable, 
                                                               m1_inst_wa, m1_inst_ra, 
                                                               m1_inst_row_repair_in, 
                                                               m1_inst_global_rrow_en_in, 
                                                               m1_inst_col_repair_in, 
                                                               m1_inst_isolation_control_in, 
                                                               m1_inst_dpslp_or_shutoffout, 
                                                               m1_inst_shutoffout, 
                                                               m1_inst_q, m2_inst_wen, 
                                                               m2_inst_ren, m2_inst_adr, 
                                                               m2_inst_din, m2_inst_async_rst, 
                                                               m2_inst_fastsleep, 
                                                               m2_inst_deepsleep, 
                                                               m2_inst_sbc, m2_inst_shutoff, 
                                                               m2_inst_mce, m2_inst_stbyp, 
                                                               m2_inst_rmce, m2_inst_wmce, 
                                                               m2_inst_wpulse, 
                                                               m2_inst_wa_disable, 
                                                               m2_inst_wa, m2_inst_ra, 
                                                               m2_inst_row_repair_in, 
                                                               m2_inst_global_rrow_en_in, 
                                                               m2_inst_col_repair_in, 
                                                               m2_inst_isolation_control_in, 
                                                               m2_inst_dpslp_or_shutoffout, 
                                                               m2_inst_shutoffout, 
                                                               m2_inst_q, m3_inst_wen, 
                                                               m3_inst_ren, m3_inst_adr, 
                                                               m3_inst_din, m3_inst_async_rst, 
                                                               m3_inst_fastsleep, 
                                                               m3_inst_deepsleep, 
                                                               m3_inst_sbc, m3_inst_shutoff, 
                                                               m3_inst_mce, m3_inst_stbyp, 
                                                               m3_inst_rmce, m3_inst_wmce, 
                                                               m3_inst_wpulse, 
                                                               m3_inst_wa_disable, 
                                                               m3_inst_wa, m3_inst_ra, 
                                                               m3_inst_row_repair_in, 
                                                               m3_inst_global_rrow_en_in, 
                                                               m3_inst_col_repair_in, 
                                                               m3_inst_isolation_control_in, 
                                                               m3_inst_dpslp_or_shutoffout, 
                                                               m3_inst_shutoffout, 
                                                               m3_inst_q, m4_inst_wen, 
                                                               m4_inst_ren, m4_inst_adr, 
                                                               m4_inst_din, m4_inst_async_rst, 
                                                               m4_inst_fastsleep, 
                                                               m4_inst_deepsleep, 
                                                               m4_inst_sbc, m4_inst_shutoff, 
                                                               m4_inst_mce, m4_inst_stbyp, 
                                                               m4_inst_rmce, m4_inst_wmce, 
                                                               m4_inst_wpulse, 
                                                               m4_inst_wa_disable, 
                                                               m4_inst_wa, m4_inst_ra, 
                                                               m4_inst_row_repair_in, 
                                                               m4_inst_global_rrow_en_in, 
                                                               m4_inst_col_repair_in, 
                                                               m4_inst_isolation_control_in, 
                                                               m4_inst_dpslp_or_shutoffout, 
                                                               m4_inst_shutoffout, 
                                                               m4_inst_q, m5_inst_wen, 
                                                               m5_inst_ren, m5_inst_adr, 
                                                               m5_inst_din, m5_inst_async_rst, 
                                                               m5_inst_fastsleep, 
                                                               m5_inst_deepsleep, 
                                                               m5_inst_sbc, m5_inst_shutoff, 
                                                               m5_inst_mce, m5_inst_stbyp, 
                                                               m5_inst_rmce, m5_inst_wmce, 
                                                               m5_inst_wpulse, 
                                                               m5_inst_wa_disable, 
                                                               m5_inst_wa, m5_inst_ra, 
                                                               m5_inst_row_repair_in, 
                                                               m5_inst_global_rrow_en_in, 
                                                               m5_inst_col_repair_in, 
                                                               m5_inst_isolation_control_in, 
                                                               m5_inst_dpslp_or_shutoffout, 
                                                               m5_inst_shutoffout, 
                                                               m5_inst_q, m6_inst_wen, 
                                                               m6_inst_ren, m6_inst_adr, 
                                                               m6_inst_din, m6_inst_async_rst, 
                                                               m6_inst_fastsleep, 
                                                               m6_inst_deepsleep, 
                                                               m6_inst_sbc, m6_inst_shutoff, 
                                                               m6_inst_mce, m6_inst_stbyp, 
                                                               m6_inst_rmce, m6_inst_wmce, 
                                                               m6_inst_wpulse, 
                                                               m6_inst_wa_disable, 
                                                               m6_inst_wa, m6_inst_ra, 
                                                               m6_inst_row_repair_in, 
                                                               m6_inst_global_rrow_en_in, 
                                                               m6_inst_col_repair_in, 
                                                               m6_inst_isolation_control_in, 
                                                               m6_inst_dpslp_or_shutoffout, 
                                                               m6_inst_shutoffout, 
                                                               m6_inst_q, m7_inst_wen, 
                                                               m7_inst_ren, m7_inst_adr, 
                                                               m7_inst_din, m7_inst_async_rst, 
                                                               m7_inst_fastsleep, 
                                                               m7_inst_deepsleep, 
                                                               m7_inst_sbc, m7_inst_shutoff, 
                                                               m7_inst_mce, m7_inst_stbyp, 
                                                               m7_inst_rmce, m7_inst_wmce, 
                                                               m7_inst_wpulse, 
                                                               m7_inst_wa_disable, 
                                                               m7_inst_wa, m7_inst_ra, 
                                                               m7_inst_row_repair_in, 
                                                               m7_inst_global_rrow_en_in, 
                                                               m7_inst_col_repair_in, 
                                                               m7_inst_isolation_control_in, 
                                                               m7_inst_dpslp_or_shutoffout, 
                                                               m7_inst_shutoffout, 
                                                               m7_inst_q, m8_inst_wen, 
                                                               m8_inst_ren, m8_inst_adr, 
                                                               m8_inst_din, m8_inst_async_rst, 
                                                               m8_inst_fastsleep, 
                                                               m8_inst_deepsleep, 
                                                               m8_inst_sbc, m8_inst_shutoff, 
                                                               m8_inst_mce, m8_inst_stbyp, 
                                                               m8_inst_rmce, m8_inst_wmce, 
                                                               m8_inst_wpulse, 
                                                               m8_inst_wa_disable, 
                                                               m8_inst_wa, m8_inst_ra, 
                                                               m8_inst_row_repair_in, 
                                                               m8_inst_global_rrow_en_in, 
                                                               m8_inst_col_repair_in, 
                                                               m8_inst_isolation_control_in, 
                                                               m8_inst_dpslp_or_shutoffout, 
                                                               m8_inst_shutoffout, 
                                                               m8_inst_q, m9_inst_wen, 
                                                               m9_inst_ren, m9_inst_adr, 
                                                               m9_inst_din, m9_inst_async_rst, 
                                                               m9_inst_fastsleep, 
                                                               m9_inst_deepsleep, 
                                                               m9_inst_sbc, m9_inst_shutoff, 
                                                               m9_inst_mce, m9_inst_stbyp, 
                                                               m9_inst_rmce, m9_inst_wmce, 
                                                               m9_inst_wpulse, 
                                                               m9_inst_wa_disable, 
                                                               m9_inst_wa, m9_inst_ra, 
                                                               m9_inst_row_repair_in, 
                                                               m9_inst_global_rrow_en_in, 
                                                               m9_inst_col_repair_in, 
                                                               m9_inst_isolation_control_in, 
                                                               m9_inst_dpslp_or_shutoffout, 
                                                               m9_inst_shutoffout, 
                                                               m9_inst_q, m10_inst_wen, 
                                                               m10_inst_ren, m10_inst_adr, 
                                                               m10_inst_din, m10_inst_async_rst, 
                                                               m10_inst_fastsleep, 
                                                               m10_inst_deepsleep, 
                                                               m10_inst_sbc, m10_inst_shutoff, 
                                                               m10_inst_mce, m10_inst_stbyp, 
                                                               m10_inst_rmce, m10_inst_wmce, 
                                                               m10_inst_wpulse, 
                                                               m10_inst_wa_disable, 
                                                               m10_inst_wa, m10_inst_ra, 
                                                               m10_inst_row_repair_in, 
                                                               m10_inst_global_rrow_en_in, 
                                                               m10_inst_col_repair_in, 
                                                               m10_inst_isolation_control_in, 
                                                               m10_inst_dpslp_or_shutoffout, 
                                                               m10_inst_shutoffout, 
                                                               m10_inst_q, m11_inst_wen, 
                                                               m11_inst_ren, m11_inst_adr, 
                                                               m11_inst_din, m11_inst_async_rst, 
                                                               m11_inst_fastsleep, 
                                                               m11_inst_deepsleep, 
                                                               m11_inst_sbc, m11_inst_shutoff, 
                                                               m11_inst_mce, m11_inst_stbyp, 
                                                               m11_inst_rmce, m11_inst_wmce, 
                                                               m11_inst_wpulse, 
                                                               m11_inst_wa_disable, 
                                                               m11_inst_wa, m11_inst_ra, 
                                                               m11_inst_row_repair_in, 
                                                               m11_inst_global_rrow_en_in, 
                                                               m11_inst_col_repair_in, 
                                                               m11_inst_isolation_control_in, 
                                                               m11_inst_dpslp_or_shutoffout, 
                                                               m11_inst_shutoffout, 
                                                               m11_inst_q, m12_inst_wen, 
                                                               m12_inst_ren, m12_inst_adr, 
                                                               m12_inst_din, m12_inst_async_rst, 
                                                               m12_inst_fastsleep, 
                                                               m12_inst_deepsleep, 
                                                               m12_inst_sbc, m12_inst_shutoff, 
                                                               m12_inst_mce, m12_inst_stbyp, 
                                                               m12_inst_rmce, m12_inst_wmce, 
                                                               m12_inst_wpulse, 
                                                               m12_inst_wa_disable, 
                                                               m12_inst_wa, m12_inst_ra, 
                                                               m12_inst_row_repair_in, 
                                                               m12_inst_global_rrow_en_in, 
                                                               m12_inst_col_repair_in, 
                                                               m12_inst_isolation_control_in, 
                                                               m12_inst_dpslp_or_shutoffout, 
                                                               m12_inst_shutoffout, 
                                                               m12_inst_q, m13_inst_wen, 
                                                               m13_inst_ren, m13_inst_adr, 
                                                               m13_inst_din, m13_inst_async_rst, 
                                                               m13_inst_fastsleep, 
                                                               m13_inst_deepsleep, 
                                                               m13_inst_sbc, m13_inst_shutoff, 
                                                               m13_inst_mce, m13_inst_stbyp, 
                                                               m13_inst_rmce, m13_inst_wmce, 
                                                               m13_inst_wpulse, 
                                                               m13_inst_wa_disable, 
                                                               m13_inst_wa, m13_inst_ra, 
                                                               m13_inst_row_repair_in, 
                                                               m13_inst_global_rrow_en_in, 
                                                               m13_inst_col_repair_in, 
                                                               m13_inst_isolation_control_in, 
                                                               m13_inst_dpslp_or_shutoffout, 
                                                               m13_inst_shutoffout, 
                                                               m13_inst_q, m14_inst_wen, 
                                                               m14_inst_ren, m14_inst_adr, 
                                                               m14_inst_din, m14_inst_async_rst, 
                                                               m14_inst_fastsleep, 
                                                               m14_inst_deepsleep, 
                                                               m14_inst_sbc, m14_inst_shutoff, 
                                                               m14_inst_mce, m14_inst_stbyp, 
                                                               m14_inst_rmce, m14_inst_wmce, 
                                                               m14_inst_wpulse, 
                                                               m14_inst_wa_disable, 
                                                               m14_inst_wa, m14_inst_ra, 
                                                               m14_inst_row_repair_in, 
                                                               m14_inst_global_rrow_en_in, 
                                                               m14_inst_col_repair_in, 
                                                               m14_inst_isolation_control_in, 
                                                               m14_inst_dpslp_or_shutoffout, 
                                                               m14_inst_shutoffout, 
                                                               m14_inst_q, m15_inst_wen, 
                                                               m15_inst_ren, m15_inst_adr, 
                                                               m15_inst_din, m15_inst_async_rst, 
                                                               m15_inst_fastsleep, 
                                                               m15_inst_deepsleep, 
                                                               m15_inst_sbc, m15_inst_shutoff, 
                                                               m15_inst_mce, m15_inst_stbyp, 
                                                               m15_inst_rmce, m15_inst_wmce, 
                                                               m15_inst_wpulse, 
                                                               m15_inst_wa_disable, 
                                                               m15_inst_wa, m15_inst_ra, 
                                                               m15_inst_row_repair_in, 
                                                               m15_inst_global_rrow_en_in, 
                                                               m15_inst_col_repair_in, 
                                                               m15_inst_isolation_control_in, 
                                                               m15_inst_dpslp_or_shutoffout, 
                                                               m15_inst_shutoffout, 
                                                               m15_inst_q, m16_inst_wen, 
                                                               m16_inst_ren, m16_inst_adr, 
                                                               m16_inst_din, m16_inst_async_rst, 
                                                               m16_inst_fastsleep, 
                                                               m16_inst_deepsleep, 
                                                               m16_inst_sbc, m16_inst_shutoff, 
                                                               m16_inst_mce, m16_inst_stbyp, 
                                                               m16_inst_rmce, m16_inst_wmce, 
                                                               m16_inst_wpulse, 
                                                               m16_inst_wa_disable, 
                                                               m16_inst_wa, m16_inst_ra, 
                                                               m16_inst_row_repair_in, 
                                                               m16_inst_global_rrow_en_in, 
                                                               m16_inst_col_repair_in, 
                                                               m16_inst_isolation_control_in, 
                                                               m16_inst_dpslp_or_shutoffout, 
                                                               m16_inst_shutoffout, 
                                                               m16_inst_q, m17_inst_wen, 
                                                               m17_inst_ren, m17_inst_adr, 
                                                               m17_inst_din, m17_inst_async_rst, 
                                                               m17_inst_fastsleep, 
                                                               m17_inst_deepsleep, 
                                                               m17_inst_sbc, m17_inst_shutoff, 
                                                               m17_inst_mce, m17_inst_stbyp, 
                                                               m17_inst_rmce, m17_inst_wmce, 
                                                               m17_inst_wpulse, 
                                                               m17_inst_wa_disable, 
                                                               m17_inst_wa, m17_inst_ra, 
                                                               m17_inst_row_repair_in, 
                                                               m17_inst_global_rrow_en_in, 
                                                               m17_inst_col_repair_in, 
                                                               m17_inst_isolation_control_in, 
                                                               m17_inst_dpslp_or_shutoffout, 
                                                               m17_inst_shutoffout, 
                                                               m17_inst_q, m18_inst_wen, 
                                                               m18_inst_ren, m18_inst_adr, 
                                                               m18_inst_din, m18_inst_async_rst, 
                                                               m18_inst_fastsleep, 
                                                               m18_inst_deepsleep, 
                                                               m18_inst_sbc, m18_inst_shutoff, 
                                                               m18_inst_mce, m18_inst_stbyp, 
                                                               m18_inst_rmce, m18_inst_wmce, 
                                                               m18_inst_wpulse, 
                                                               m18_inst_wa_disable, 
                                                               m18_inst_wa, m18_inst_ra, 
                                                               m18_inst_row_repair_in, 
                                                               m18_inst_global_rrow_en_in, 
                                                               m18_inst_col_repair_in, 
                                                               m18_inst_isolation_control_in, 
                                                               m18_inst_dpslp_or_shutoffout, 
                                                               m18_inst_shutoffout, 
                                                               m18_inst_q, m19_inst_wen, 
                                                               m19_inst_ren, m19_inst_adr, 
                                                               m19_inst_din, m19_inst_async_rst, 
                                                               m19_inst_fastsleep, 
                                                               m19_inst_deepsleep, 
                                                               m19_inst_sbc, m19_inst_shutoff, 
                                                               m19_inst_mce, m19_inst_stbyp, 
                                                               m19_inst_rmce, m19_inst_wmce, 
                                                               m19_inst_wpulse, 
                                                               m19_inst_wa_disable, 
                                                               m19_inst_wa, m19_inst_ra, 
                                                               m19_inst_row_repair_in, 
                                                               m19_inst_global_rrow_en_in, 
                                                               m19_inst_col_repair_in, 
                                                               m19_inst_isolation_control_in, 
                                                               m19_inst_dpslp_or_shutoffout, 
                                                               m19_inst_shutoffout, 
                                                               m19_inst_q, m20_inst_wen, 
                                                               m20_inst_ren, m20_inst_adr, 
                                                               m20_inst_din, m20_inst_async_rst, 
                                                               m20_inst_fastsleep, 
                                                               m20_inst_deepsleep, 
                                                               m20_inst_sbc, m20_inst_shutoff, 
                                                               m20_inst_mce, m20_inst_stbyp, 
                                                               m20_inst_rmce, m20_inst_wmce, 
                                                               m20_inst_wpulse, 
                                                               m20_inst_wa_disable, 
                                                               m20_inst_wa, m20_inst_ra, 
                                                               m20_inst_row_repair_in, 
                                                               m20_inst_global_rrow_en_in, 
                                                               m20_inst_col_repair_in, 
                                                               m20_inst_isolation_control_in, 
                                                               m20_inst_dpslp_or_shutoffout, 
                                                               m20_inst_shutoffout, 
                                                               m20_inst_q, m21_inst_wen, 
                                                               m21_inst_ren, m21_inst_adr, 
                                                               m21_inst_din, m21_inst_async_rst, 
                                                               m21_inst_fastsleep, 
                                                               m21_inst_deepsleep, 
                                                               m21_inst_sbc, m21_inst_shutoff, 
                                                               m21_inst_mce, m21_inst_stbyp, 
                                                               m21_inst_rmce, m21_inst_wmce, 
                                                               m21_inst_wpulse, 
                                                               m21_inst_wa_disable, 
                                                               m21_inst_wa, m21_inst_ra, 
                                                               m21_inst_row_repair_in, 
                                                               m21_inst_global_rrow_en_in, 
                                                               m21_inst_col_repair_in, 
                                                               m21_inst_isolation_control_in, 
                                                               m21_inst_dpslp_or_shutoffout, 
                                                               m21_inst_shutoffout, 
                                                               m21_inst_q, m22_inst_wen, 
                                                               m22_inst_ren, m22_inst_adr, 
                                                               m22_inst_din, m22_inst_async_rst, 
                                                               m22_inst_fastsleep, 
                                                               m22_inst_deepsleep, 
                                                               m22_inst_sbc, m22_inst_shutoff, 
                                                               m22_inst_mce, m22_inst_stbyp, 
                                                               m22_inst_rmce, m22_inst_wmce, 
                                                               m22_inst_wpulse, 
                                                               m22_inst_wa_disable, 
                                                               m22_inst_wa, m22_inst_ra, 
                                                               m22_inst_row_repair_in, 
                                                               m22_inst_global_rrow_en_in, 
                                                               m22_inst_col_repair_in, 
                                                               m22_inst_isolation_control_in, 
                                                               m22_inst_dpslp_or_shutoffout, 
                                                               m22_inst_shutoffout, 
                                                               m22_inst_q, m23_inst_wen, 
                                                               m23_inst_ren, m23_inst_adr, 
                                                               m23_inst_din, m23_inst_async_rst, 
                                                               m23_inst_fastsleep, 
                                                               m23_inst_deepsleep, 
                                                               m23_inst_sbc, m23_inst_shutoff, 
                                                               m23_inst_mce, m23_inst_stbyp, 
                                                               m23_inst_rmce, m23_inst_wmce, 
                                                               m23_inst_wpulse, 
                                                               m23_inst_wa_disable, 
                                                               m23_inst_wa, m23_inst_ra, 
                                                               m23_inst_row_repair_in, 
                                                               m23_inst_global_rrow_en_in, 
                                                               m23_inst_col_repair_in, 
                                                               m23_inst_isolation_control_in, 
                                                               m23_inst_dpslp_or_shutoffout, 
                                                               m23_inst_shutoffout, 
                                                               m23_inst_q, m24_inst_wen, 
                                                               m24_inst_ren, m24_inst_adr, 
                                                               m24_inst_din, m24_inst_async_rst, 
                                                               m24_inst_fastsleep, 
                                                               m24_inst_deepsleep, 
                                                               m24_inst_sbc, m24_inst_shutoff, 
                                                               m24_inst_mce, m24_inst_stbyp, 
                                                               m24_inst_rmce, m24_inst_wmce, 
                                                               m24_inst_wpulse, 
                                                               m24_inst_wa_disable, 
                                                               m24_inst_wa, m24_inst_ra, 
                                                               m24_inst_row_repair_in, 
                                                               m24_inst_global_rrow_en_in, 
                                                               m24_inst_col_repair_in, 
                                                               m24_inst_isolation_control_in, 
                                                               m24_inst_dpslp_or_shutoffout, 
                                                               m24_inst_shutoffout, 
                                                               m24_inst_q, m25_inst_wen, 
                                                               m25_inst_ren, m25_inst_adr, 
                                                               m25_inst_din, m25_inst_async_rst, 
                                                               m25_inst_fastsleep, 
                                                               m25_inst_deepsleep, 
                                                               m25_inst_sbc, m25_inst_shutoff, 
                                                               m25_inst_mce, m25_inst_stbyp, 
                                                               m25_inst_rmce, m25_inst_wmce, 
                                                               m25_inst_wpulse, 
                                                               m25_inst_wa_disable, 
                                                               m25_inst_wa, m25_inst_ra, 
                                                               m25_inst_row_repair_in, 
                                                               m25_inst_global_rrow_en_in, 
                                                               m25_inst_col_repair_in, 
                                                               m25_inst_isolation_control_in, 
                                                               m25_inst_dpslp_or_shutoffout, 
                                                               m25_inst_shutoffout, 
                                                               m25_inst_q, m26_inst_wen, 
                                                               m26_inst_ren, m26_inst_adr, 
                                                               m26_inst_din, m26_inst_async_rst, 
                                                               m26_inst_fastsleep, 
                                                               m26_inst_deepsleep, 
                                                               m26_inst_sbc, m26_inst_shutoff, 
                                                               m26_inst_mce, m26_inst_stbyp, 
                                                               m26_inst_rmce, m26_inst_wmce, 
                                                               m26_inst_wpulse, 
                                                               m26_inst_wa_disable, 
                                                               m26_inst_wa, m26_inst_ra, 
                                                               m26_inst_row_repair_in, 
                                                               m26_inst_global_rrow_en_in, 
                                                               m26_inst_col_repair_in, 
                                                               m26_inst_isolation_control_in, 
                                                               m26_inst_dpslp_or_shutoffout, 
                                                               m26_inst_shutoffout, 
                                                               m26_inst_q, m27_inst_wen, 
                                                               m27_inst_ren, m27_inst_adr, 
                                                               m27_inst_din, m27_inst_async_rst, 
                                                               m27_inst_fastsleep, 
                                                               m27_inst_deepsleep, 
                                                               m27_inst_sbc, m27_inst_shutoff, 
                                                               m27_inst_mce, m27_inst_stbyp, 
                                                               m27_inst_rmce, m27_inst_wmce, 
                                                               m27_inst_wpulse, 
                                                               m27_inst_wa_disable, 
                                                               m27_inst_wa, m27_inst_ra, 
                                                               m27_inst_row_repair_in, 
                                                               m27_inst_global_rrow_en_in, 
                                                               m27_inst_col_repair_in, 
                                                               m27_inst_isolation_control_in, 
                                                               m27_inst_dpslp_or_shutoffout, 
                                                               m27_inst_shutoffout, 
                                                               m27_inst_q, m28_inst_wen, 
                                                               m28_inst_ren, m28_inst_adr, 
                                                               m28_inst_din, m28_inst_async_rst, 
                                                               m28_inst_fastsleep, 
                                                               m28_inst_deepsleep, 
                                                               m28_inst_sbc, m28_inst_shutoff, 
                                                               m28_inst_mce, m28_inst_stbyp, 
                                                               m28_inst_rmce, m28_inst_wmce, 
                                                               m28_inst_wpulse, 
                                                               m28_inst_wa_disable, 
                                                               m28_inst_wa, m28_inst_ra, 
                                                               m28_inst_row_repair_in, 
                                                               m28_inst_global_rrow_en_in, 
                                                               m28_inst_col_repair_in, 
                                                               m28_inst_isolation_control_in, 
                                                               m28_inst_dpslp_or_shutoffout, 
                                                               m28_inst_shutoffout, 
                                                               m28_inst_q, m29_inst_wen, 
                                                               m29_inst_ren, m29_inst_adr, 
                                                               m29_inst_din, m29_inst_async_rst, 
                                                               m29_inst_fastsleep, 
                                                               m29_inst_deepsleep, 
                                                               m29_inst_sbc, m29_inst_shutoff, 
                                                               m29_inst_mce, m29_inst_stbyp, 
                                                               m29_inst_rmce, m29_inst_wmce, 
                                                               m29_inst_wpulse, 
                                                               m29_inst_wa_disable, 
                                                               m29_inst_wa, m29_inst_ra, 
                                                               m29_inst_row_repair_in, 
                                                               m29_inst_global_rrow_en_in, 
                                                               m29_inst_col_repair_in, 
                                                               m29_inst_isolation_control_in, 
                                                               m29_inst_dpslp_or_shutoffout, 
                                                               m29_inst_shutoffout, 
                                                               m29_inst_q, m30_inst_wen, 
                                                               m30_inst_ren, m30_inst_adr, 
                                                               m30_inst_din, m30_inst_async_rst, 
                                                               m30_inst_fastsleep, 
                                                               m30_inst_deepsleep, 
                                                               m30_inst_sbc, m30_inst_shutoff, 
                                                               m30_inst_mce, m30_inst_stbyp, 
                                                               m30_inst_rmce, m30_inst_wmce, 
                                                               m30_inst_wpulse, 
                                                               m30_inst_wa_disable, 
                                                               m30_inst_wa, m30_inst_ra, 
                                                               m30_inst_row_repair_in, 
                                                               m30_inst_global_rrow_en_in, 
                                                               m30_inst_col_repair_in, 
                                                               m30_inst_isolation_control_in, 
                                                               m30_inst_dpslp_or_shutoffout, 
                                                               m30_inst_shutoffout, 
                                                               m30_inst_q, m31_inst_wen, 
                                                               m31_inst_ren, m31_inst_adr, 
                                                               m31_inst_din, m31_inst_async_rst, 
                                                               m31_inst_fastsleep, 
                                                               m31_inst_deepsleep, 
                                                               m31_inst_sbc, m31_inst_shutoff, 
                                                               m31_inst_mce, m31_inst_stbyp, 
                                                               m31_inst_rmce, m31_inst_wmce, 
                                                               m31_inst_wpulse, 
                                                               m31_inst_wa_disable, 
                                                               m31_inst_wa, m31_inst_ra, 
                                                               m31_inst_row_repair_in, 
                                                               m31_inst_global_rrow_en_in, 
                                                               m31_inst_col_repair_in, 
                                                               m31_inst_isolation_control_in, 
                                                               m31_inst_dpslp_or_shutoffout, 
                                                               m31_inst_shutoffout, 
                                                               m31_inst_q, m32_inst_wen, 
                                                               m32_inst_ren, m32_inst_adr, 
                                                               m32_inst_din, m32_inst_async_rst, 
                                                               m32_inst_fastsleep, 
                                                               m32_inst_deepsleep, 
                                                               m32_inst_sbc, m32_inst_shutoff, 
                                                               m32_inst_mce, m32_inst_stbyp, 
                                                               m32_inst_rmce, m32_inst_wmce, 
                                                               m32_inst_wpulse, 
                                                               m32_inst_wa_disable, 
                                                               m32_inst_wa, m32_inst_ra, 
                                                               m32_inst_row_repair_in, 
                                                               m32_inst_global_rrow_en_in, 
                                                               m32_inst_col_repair_in, 
                                                               m32_inst_isolation_control_in, 
                                                               m32_inst_dpslp_or_shutoffout, 
                                                               m32_inst_shutoffout, 
                                                               m32_inst_q, m33_inst_wen, 
                                                               m33_inst_ren, m33_inst_adr, 
                                                               m33_inst_din, m33_inst_async_rst, 
                                                               m33_inst_fastsleep, 
                                                               m33_inst_deepsleep, 
                                                               m33_inst_sbc, m33_inst_shutoff, 
                                                               m33_inst_mce, m33_inst_stbyp, 
                                                               m33_inst_rmce, m33_inst_wmce, 
                                                               m33_inst_wpulse, 
                                                               m33_inst_wa_disable, 
                                                               m33_inst_wa, m33_inst_ra, 
                                                               m33_inst_row_repair_in, 
                                                               m33_inst_global_rrow_en_in, 
                                                               m33_inst_col_repair_in, 
                                                               m33_inst_isolation_control_in, 
                                                               m33_inst_dpslp_or_shutoffout, 
                                                               m33_inst_shutoffout, 
                                                               m33_inst_q, m34_inst_wen, 
                                                               m34_inst_ren, m34_inst_adr, 
                                                               m34_inst_din, m34_inst_async_rst, 
                                                               m34_inst_fastsleep, 
                                                               m34_inst_deepsleep, 
                                                               m34_inst_sbc, m34_inst_shutoff, 
                                                               m34_inst_mce, m34_inst_stbyp, 
                                                               m34_inst_rmce, m34_inst_wmce, 
                                                               m34_inst_wpulse, 
                                                               m34_inst_wa_disable, 
                                                               m34_inst_wa, m34_inst_ra, 
                                                               m34_inst_row_repair_in, 
                                                               m34_inst_global_rrow_en_in, 
                                                               m34_inst_col_repair_in, 
                                                               m34_inst_isolation_control_in, 
                                                               m34_inst_dpslp_or_shutoffout, 
                                                               m34_inst_shutoffout, 
                                                               m34_inst_q, m35_inst_wen, 
                                                               m35_inst_ren, m35_inst_adr, 
                                                               m35_inst_din, m35_inst_async_rst, 
                                                               m35_inst_fastsleep, 
                                                               m35_inst_deepsleep, 
                                                               m35_inst_sbc, m35_inst_shutoff, 
                                                               m35_inst_mce, m35_inst_stbyp, 
                                                               m35_inst_rmce, m35_inst_wmce, 
                                                               m35_inst_wpulse, 
                                                               m35_inst_wa_disable, 
                                                               m35_inst_wa, m35_inst_ra, 
                                                               m35_inst_row_repair_in, 
                                                               m35_inst_global_rrow_en_in, 
                                                               m35_inst_col_repair_in, 
                                                               m35_inst_isolation_control_in, 
                                                               m35_inst_dpslp_or_shutoffout, 
                                                               m35_inst_shutoffout, 
                                                               m35_inst_q, m36_inst_wen, 
                                                               m36_inst_ren, m36_inst_adr, 
                                                               m36_inst_din, m36_inst_async_rst, 
                                                               m36_inst_fastsleep, 
                                                               m36_inst_deepsleep, 
                                                               m36_inst_sbc, m36_inst_shutoff, 
                                                               m36_inst_mce, m36_inst_stbyp, 
                                                               m36_inst_rmce, m36_inst_wmce, 
                                                               m36_inst_wpulse, 
                                                               m36_inst_wa_disable, 
                                                               m36_inst_wa, m36_inst_ra, 
                                                               m36_inst_row_repair_in, 
                                                               m36_inst_global_rrow_en_in, 
                                                               m36_inst_col_repair_in, 
                                                               m36_inst_isolation_control_in, 
                                                               m36_inst_dpslp_or_shutoffout, 
                                                               m36_inst_shutoffout, 
                                                               m36_inst_q, m37_inst_wen, 
                                                               m37_inst_ren, m37_inst_adr, 
                                                               m37_inst_din, m37_inst_async_rst, 
                                                               m37_inst_fastsleep, 
                                                               m37_inst_deepsleep, 
                                                               m37_inst_sbc, m37_inst_shutoff, 
                                                               m37_inst_mce, m37_inst_stbyp, 
                                                               m37_inst_rmce, m37_inst_wmce, 
                                                               m37_inst_wpulse, 
                                                               m37_inst_wa_disable, 
                                                               m37_inst_wa, m37_inst_ra, 
                                                               m37_inst_row_repair_in, 
                                                               m37_inst_global_rrow_en_in, 
                                                               m37_inst_col_repair_in, 
                                                               m37_inst_isolation_control_in, 
                                                               m37_inst_dpslp_or_shutoffout, 
                                                               m37_inst_shutoffout, 
                                                               m37_inst_q, m38_inst_wen, 
                                                               m38_inst_ren, m38_inst_adr, 
                                                               m38_inst_din, m38_inst_async_rst, 
                                                               m38_inst_fastsleep, 
                                                               m38_inst_deepsleep, 
                                                               m38_inst_sbc, m38_inst_shutoff, 
                                                               m38_inst_mce, m38_inst_stbyp, 
                                                               m38_inst_rmce, m38_inst_wmce, 
                                                               m38_inst_wpulse, 
                                                               m38_inst_wa_disable, 
                                                               m38_inst_wa, m38_inst_ra, 
                                                               m38_inst_row_repair_in, 
                                                               m38_inst_global_rrow_en_in, 
                                                               m38_inst_col_repair_in, 
                                                               m38_inst_isolation_control_in, 
                                                               m38_inst_dpslp_or_shutoffout, 
                                                               m38_inst_shutoffout, 
                                                               m38_inst_q, m39_inst_wen, 
                                                               m39_inst_ren, m39_inst_adr, 
                                                               m39_inst_din, m39_inst_async_rst, 
                                                               m39_inst_fastsleep, 
                                                               m39_inst_deepsleep, 
                                                               m39_inst_sbc, m39_inst_shutoff, 
                                                               m39_inst_mce, m39_inst_stbyp, 
                                                               m39_inst_rmce, m39_inst_wmce, 
                                                               m39_inst_wpulse, 
                                                               m39_inst_wa_disable, 
                                                               m39_inst_wa, m39_inst_ra, 
                                                               m39_inst_row_repair_in, 
                                                               m39_inst_global_rrow_en_in, 
                                                               m39_inst_col_repair_in, 
                                                               m39_inst_isolation_control_in, 
                                                               m39_inst_dpslp_or_shutoffout, 
                                                               m39_inst_shutoffout, 
                                                               m39_inst_q, m40_inst_wen, 
                                                               m40_inst_ren, m40_inst_adr, 
                                                               m40_inst_din, m40_inst_async_rst, 
                                                               m40_inst_fastsleep, 
                                                               m40_inst_deepsleep, 
                                                               m40_inst_sbc, m40_inst_shutoff, 
                                                               m40_inst_mce, m40_inst_stbyp, 
                                                               m40_inst_rmce, m40_inst_wmce, 
                                                               m40_inst_wpulse, 
                                                               m40_inst_wa_disable, 
                                                               m40_inst_wa, m40_inst_ra, 
                                                               m40_inst_row_repair_in, 
                                                               m40_inst_global_rrow_en_in, 
                                                               m40_inst_col_repair_in, 
                                                               m40_inst_isolation_control_in, 
                                                               m40_inst_dpslp_or_shutoffout, 
                                                               m40_inst_shutoffout, 
                                                               m40_inst_q, reset, 
                                                               ijtag_select, si, 
                                                               capture_en, shift_en, 
                                                               update_en, tck, 
                                                               so, bisr_so, bisr_si, 
                                                               bisr_se, bisr_clock, 
                                                               bisr_clear);
  input  [71:0] m33_inst_din, m34_inst_din, m35_inst_din, m36_inst_din;
  input  [31:0] m37_inst_din, m38_inst_din, m39_inst_din, m40_inst_din;
  input  [25:0] m1_inst_row_repair_in, m2_inst_row_repair_in, 
                m3_inst_row_repair_in, m4_inst_row_repair_in, 
                m5_inst_row_repair_in, m6_inst_row_repair_in, 
                m7_inst_row_repair_in, m8_inst_row_repair_in, 
                m9_inst_row_repair_in, m10_inst_row_repair_in, 
                m11_inst_row_repair_in, m12_inst_row_repair_in, 
                m13_inst_row_repair_in, m14_inst_row_repair_in, 
                m15_inst_row_repair_in, m16_inst_row_repair_in, 
                m17_inst_row_repair_in, m18_inst_row_repair_in, 
                m19_inst_row_repair_in, m20_inst_row_repair_in, 
                m21_inst_row_repair_in, m22_inst_row_repair_in, 
                m23_inst_row_repair_in, m24_inst_row_repair_in, 
                m25_inst_row_repair_in, m26_inst_row_repair_in, 
                m27_inst_row_repair_in, m28_inst_row_repair_in, 
                m29_inst_row_repair_in, m30_inst_row_repair_in, 
                m31_inst_row_repair_in, m32_inst_row_repair_in, 
                m33_inst_row_repair_in, m34_inst_row_repair_in, 
                m35_inst_row_repair_in, m36_inst_row_repair_in, 
                m37_inst_row_repair_in, m38_inst_row_repair_in, 
                m39_inst_row_repair_in, m40_inst_row_repair_in;
  input  [21:0] m1_inst_din, m2_inst_din, m3_inst_din, m4_inst_din, 
                m5_inst_din, m6_inst_din, m7_inst_din, m8_inst_din, 
                m9_inst_din, m10_inst_din, m11_inst_din, m12_inst_din, 
                m13_inst_din, m14_inst_din, m15_inst_din, m16_inst_din, 
                m17_inst_din, m18_inst_din, m19_inst_din, m20_inst_din, 
                m21_inst_din, m22_inst_din, m23_inst_din, m24_inst_din, 
                m25_inst_din, m26_inst_din, m27_inst_din, m28_inst_din, 
                m29_inst_din, m30_inst_din, m31_inst_din, m32_inst_din;
  input  [12:0] m1_inst_col_repair_in, m2_inst_col_repair_in, 
                m3_inst_col_repair_in, m4_inst_col_repair_in, 
                m5_inst_col_repair_in, m6_inst_col_repair_in, 
                m7_inst_col_repair_in, m8_inst_col_repair_in, 
                m9_inst_col_repair_in, m10_inst_col_repair_in, 
                m11_inst_col_repair_in, m12_inst_col_repair_in, 
                m13_inst_col_repair_in, m14_inst_col_repair_in, 
                m15_inst_col_repair_in, m16_inst_col_repair_in, 
                m17_inst_col_repair_in, m18_inst_col_repair_in, 
                m19_inst_col_repair_in, m20_inst_col_repair_in, 
                m21_inst_col_repair_in, m22_inst_col_repair_in, 
                m23_inst_col_repair_in, m24_inst_col_repair_in, 
                m25_inst_col_repair_in, m26_inst_col_repair_in, 
                m27_inst_col_repair_in, m28_inst_col_repair_in, 
                m29_inst_col_repair_in, m30_inst_col_repair_in, 
                m31_inst_col_repair_in, m32_inst_col_repair_in, 
                m33_inst_col_repair_in, m34_inst_col_repair_in, 
                m35_inst_col_repair_in, m36_inst_col_repair_in, 
                m37_inst_col_repair_in, m38_inst_col_repair_in, 
                m39_inst_col_repair_in, m40_inst_col_repair_in;
  input  [9:0] m1_inst_adr, m2_inst_adr, m3_inst_adr, m4_inst_adr, m5_inst_adr, 
               m6_inst_adr, m7_inst_adr, m8_inst_adr, m9_inst_adr, 
               m10_inst_adr, m11_inst_adr, m12_inst_adr, m13_inst_adr, 
               m14_inst_adr, m15_inst_adr, m16_inst_adr, m17_inst_adr, 
               m18_inst_adr, m19_inst_adr, m20_inst_adr, m21_inst_adr, 
               m22_inst_adr, m23_inst_adr, m24_inst_adr, m25_inst_adr, 
               m26_inst_adr, m27_inst_adr, m28_inst_adr, m29_inst_adr, 
               m30_inst_adr, m31_inst_adr, m32_inst_adr, m33_inst_adr, 
               m34_inst_adr, m35_inst_adr, m36_inst_adr;
  input  [8:0] m37_inst_adr, m38_inst_adr, m39_inst_adr, m40_inst_adr;
  input  [3:0] m1_inst_rmce, m2_inst_rmce, m3_inst_rmce, m4_inst_rmce, 
               m5_inst_rmce, m6_inst_rmce, m7_inst_rmce, m8_inst_rmce, 
               m9_inst_rmce, m10_inst_rmce, m11_inst_rmce, m12_inst_rmce, 
               m13_inst_rmce, m14_inst_rmce, m15_inst_rmce, m16_inst_rmce, 
               m17_inst_rmce, m18_inst_rmce, m19_inst_rmce, m20_inst_rmce, 
               m21_inst_rmce, m22_inst_rmce, m23_inst_rmce, m24_inst_rmce, 
               m25_inst_rmce, m26_inst_rmce, m27_inst_rmce, m28_inst_rmce, 
               m29_inst_rmce, m30_inst_rmce, m31_inst_rmce, m32_inst_rmce, 
               m33_inst_rmce, m34_inst_rmce, m35_inst_rmce, m36_inst_rmce, 
               m37_inst_rmce, m38_inst_rmce, m39_inst_rmce, m40_inst_rmce;
  input  [2:0] m1_inst_wa, m2_inst_wa, m3_inst_wa, m4_inst_wa, m5_inst_wa, 
               m6_inst_wa, m7_inst_wa, m8_inst_wa, m9_inst_wa, m10_inst_wa, 
               m11_inst_wa, m12_inst_wa, m13_inst_wa, m14_inst_wa, m15_inst_wa, 
               m16_inst_wa, m17_inst_wa, m18_inst_wa, m19_inst_wa, m20_inst_wa, 
               m21_inst_wa, m22_inst_wa, m23_inst_wa, m24_inst_wa, m25_inst_wa, 
               m26_inst_wa, m27_inst_wa, m28_inst_wa, m29_inst_wa, m30_inst_wa, 
               m31_inst_wa, m32_inst_wa, m33_inst_wa, m34_inst_wa, m35_inst_wa, 
               m36_inst_wa, m37_inst_wa, m38_inst_wa, m39_inst_wa, m40_inst_wa;
  input  [1:0] m1_inst_sbc, m1_inst_wmce, m1_inst_wpulse, m1_inst_ra, 
               m1_inst_global_rrow_en_in, m2_inst_sbc, m2_inst_wmce, 
               m2_inst_wpulse, m2_inst_ra, m2_inst_global_rrow_en_in, 
               m3_inst_sbc, m3_inst_wmce, m3_inst_wpulse, m3_inst_ra, 
               m3_inst_global_rrow_en_in, m4_inst_sbc, m4_inst_wmce, 
               m4_inst_wpulse, m4_inst_ra, m4_inst_global_rrow_en_in, 
               m5_inst_sbc, m5_inst_wmce, m5_inst_wpulse, m5_inst_ra, 
               m5_inst_global_rrow_en_in, m6_inst_sbc, m6_inst_wmce, 
               m6_inst_wpulse, m6_inst_ra, m6_inst_global_rrow_en_in, 
               m7_inst_sbc, m7_inst_wmce, m7_inst_wpulse, m7_inst_ra, 
               m7_inst_global_rrow_en_in, m8_inst_sbc, m8_inst_wmce, 
               m8_inst_wpulse, m8_inst_ra, m8_inst_global_rrow_en_in, 
               m9_inst_sbc, m9_inst_wmce, m9_inst_wpulse, m9_inst_ra, 
               m9_inst_global_rrow_en_in, m10_inst_sbc, m10_inst_wmce, 
               m10_inst_wpulse, m10_inst_ra, m10_inst_global_rrow_en_in, 
               m11_inst_sbc, m11_inst_wmce, m11_inst_wpulse, m11_inst_ra, 
               m11_inst_global_rrow_en_in, m12_inst_sbc, m12_inst_wmce, 
               m12_inst_wpulse, m12_inst_ra, m12_inst_global_rrow_en_in, 
               m13_inst_sbc, m13_inst_wmce, m13_inst_wpulse, m13_inst_ra, 
               m13_inst_global_rrow_en_in, m14_inst_sbc, m14_inst_wmce, 
               m14_inst_wpulse, m14_inst_ra, m14_inst_global_rrow_en_in, 
               m15_inst_sbc, m15_inst_wmce, m15_inst_wpulse, m15_inst_ra, 
               m15_inst_global_rrow_en_in, m16_inst_sbc, m16_inst_wmce, 
               m16_inst_wpulse, m16_inst_ra, m16_inst_global_rrow_en_in, 
               m17_inst_sbc, m17_inst_wmce, m17_inst_wpulse, m17_inst_ra, 
               m17_inst_global_rrow_en_in, m18_inst_sbc, m18_inst_wmce, 
               m18_inst_wpulse, m18_inst_ra, m18_inst_global_rrow_en_in, 
               m19_inst_sbc, m19_inst_wmce, m19_inst_wpulse, m19_inst_ra, 
               m19_inst_global_rrow_en_in, m20_inst_sbc, m20_inst_wmce, 
               m20_inst_wpulse, m20_inst_ra, m20_inst_global_rrow_en_in, 
               m21_inst_sbc, m21_inst_wmce, m21_inst_wpulse, m21_inst_ra, 
               m21_inst_global_rrow_en_in, m22_inst_sbc, m22_inst_wmce, 
               m22_inst_wpulse, m22_inst_ra, m22_inst_global_rrow_en_in, 
               m23_inst_sbc, m23_inst_wmce, m23_inst_wpulse, m23_inst_ra, 
               m23_inst_global_rrow_en_in, m24_inst_sbc, m24_inst_wmce, 
               m24_inst_wpulse, m24_inst_ra, m24_inst_global_rrow_en_in, 
               m25_inst_sbc, m25_inst_wmce, m25_inst_wpulse, m25_inst_ra, 
               m25_inst_global_rrow_en_in, m26_inst_sbc, m26_inst_wmce, 
               m26_inst_wpulse, m26_inst_ra, m26_inst_global_rrow_en_in, 
               m27_inst_sbc, m27_inst_wmce, m27_inst_wpulse, m27_inst_ra, 
               m27_inst_global_rrow_en_in, m28_inst_sbc, m28_inst_wmce, 
               m28_inst_wpulse, m28_inst_ra, m28_inst_global_rrow_en_in, 
               m29_inst_sbc, m29_inst_wmce, m29_inst_wpulse, m29_inst_ra, 
               m29_inst_global_rrow_en_in, m30_inst_sbc, m30_inst_wmce, 
               m30_inst_wpulse, m30_inst_ra, m30_inst_global_rrow_en_in, 
               m31_inst_sbc, m31_inst_wmce, m31_inst_wpulse, m31_inst_ra, 
               m31_inst_global_rrow_en_in, m32_inst_sbc, m32_inst_wmce, 
               m32_inst_wpulse, m32_inst_ra, m32_inst_global_rrow_en_in, 
               m33_inst_sbc, m33_inst_wmce, m33_inst_wpulse, m33_inst_ra, 
               m33_inst_global_rrow_en_in, m34_inst_sbc, m34_inst_wmce, 
               m34_inst_wpulse, m34_inst_ra, m34_inst_global_rrow_en_in, 
               m35_inst_sbc, m35_inst_wmce, m35_inst_wpulse, m35_inst_ra, 
               m35_inst_global_rrow_en_in, m36_inst_sbc, m36_inst_wmce, 
               m36_inst_wpulse, m36_inst_ra, m36_inst_global_rrow_en_in, 
               m37_inst_sbc, m37_inst_wmce, m37_inst_wpulse, m37_inst_ra, 
               m37_inst_global_rrow_en_in, m38_inst_sbc, m38_inst_wmce, 
               m38_inst_wpulse, m38_inst_ra, m38_inst_global_rrow_en_in, 
               m39_inst_sbc, m39_inst_wmce, m39_inst_wpulse, m39_inst_ra, 
               m39_inst_global_rrow_en_in, m40_inst_sbc, m40_inst_wmce, 
               m40_inst_wpulse, m40_inst_ra, m40_inst_global_rrow_en_in;
  input  LV_TM, MEM_BYPASS_EN, SCAN_SHIFT_EN, MCP_BOUNDING_EN, clk_clk_bbm, 
         m1_inst_wen, m1_inst_ren, m1_inst_async_rst, m1_inst_fastsleep, 
         m1_inst_deepsleep, m1_inst_shutoff, m1_inst_mce, m1_inst_stbyp, 
         m1_inst_wa_disable, m1_inst_isolation_control_in, m2_inst_wen, 
         m2_inst_ren, m2_inst_async_rst, m2_inst_fastsleep, m2_inst_deepsleep, 
         m2_inst_shutoff, m2_inst_mce, m2_inst_stbyp, m2_inst_wa_disable, 
         m2_inst_isolation_control_in, m3_inst_wen, m3_inst_ren, 
         m3_inst_async_rst, m3_inst_fastsleep, m3_inst_deepsleep, 
         m3_inst_shutoff, m3_inst_mce, m3_inst_stbyp, m3_inst_wa_disable, 
         m3_inst_isolation_control_in, m4_inst_wen, m4_inst_ren, 
         m4_inst_async_rst, m4_inst_fastsleep, m4_inst_deepsleep, 
         m4_inst_shutoff, m4_inst_mce, m4_inst_stbyp, m4_inst_wa_disable, 
         m4_inst_isolation_control_in, m5_inst_wen, m5_inst_ren, 
         m5_inst_async_rst, m5_inst_fastsleep, m5_inst_deepsleep, 
         m5_inst_shutoff, m5_inst_mce, m5_inst_stbyp, m5_inst_wa_disable, 
         m5_inst_isolation_control_in, m6_inst_wen, m6_inst_ren, 
         m6_inst_async_rst, m6_inst_fastsleep, m6_inst_deepsleep, 
         m6_inst_shutoff, m6_inst_mce, m6_inst_stbyp, m6_inst_wa_disable, 
         m6_inst_isolation_control_in, m7_inst_wen, m7_inst_ren, 
         m7_inst_async_rst, m7_inst_fastsleep, m7_inst_deepsleep, 
         m7_inst_shutoff, m7_inst_mce, m7_inst_stbyp, m7_inst_wa_disable, 
         m7_inst_isolation_control_in, m8_inst_wen, m8_inst_ren, 
         m8_inst_async_rst, m8_inst_fastsleep, m8_inst_deepsleep, 
         m8_inst_shutoff, m8_inst_mce, m8_inst_stbyp, m8_inst_wa_disable, 
         m8_inst_isolation_control_in, m9_inst_wen, m9_inst_ren, 
         m9_inst_async_rst, m9_inst_fastsleep, m9_inst_deepsleep, 
         m9_inst_shutoff, m9_inst_mce, m9_inst_stbyp, m9_inst_wa_disable, 
         m9_inst_isolation_control_in, m10_inst_wen, m10_inst_ren, 
         m10_inst_async_rst, m10_inst_fastsleep, m10_inst_deepsleep, 
         m10_inst_shutoff, m10_inst_mce, m10_inst_stbyp, m10_inst_wa_disable, 
         m10_inst_isolation_control_in, m11_inst_wen, m11_inst_ren, 
         m11_inst_async_rst, m11_inst_fastsleep, m11_inst_deepsleep, 
         m11_inst_shutoff, m11_inst_mce, m11_inst_stbyp, m11_inst_wa_disable, 
         m11_inst_isolation_control_in, m12_inst_wen, m12_inst_ren, 
         m12_inst_async_rst, m12_inst_fastsleep, m12_inst_deepsleep, 
         m12_inst_shutoff, m12_inst_mce, m12_inst_stbyp, m12_inst_wa_disable, 
         m12_inst_isolation_control_in, m13_inst_wen, m13_inst_ren, 
         m13_inst_async_rst, m13_inst_fastsleep, m13_inst_deepsleep, 
         m13_inst_shutoff, m13_inst_mce, m13_inst_stbyp, m13_inst_wa_disable, 
         m13_inst_isolation_control_in, m14_inst_wen, m14_inst_ren, 
         m14_inst_async_rst, m14_inst_fastsleep, m14_inst_deepsleep, 
         m14_inst_shutoff, m14_inst_mce, m14_inst_stbyp, m14_inst_wa_disable, 
         m14_inst_isolation_control_in, m15_inst_wen, m15_inst_ren, 
         m15_inst_async_rst, m15_inst_fastsleep, m15_inst_deepsleep, 
         m15_inst_shutoff, m15_inst_mce, m15_inst_stbyp, m15_inst_wa_disable, 
         m15_inst_isolation_control_in, m16_inst_wen, m16_inst_ren, 
         m16_inst_async_rst, m16_inst_fastsleep, m16_inst_deepsleep, 
         m16_inst_shutoff, m16_inst_mce, m16_inst_stbyp, m16_inst_wa_disable, 
         m16_inst_isolation_control_in, m17_inst_wen, m17_inst_ren, 
         m17_inst_async_rst, m17_inst_fastsleep, m17_inst_deepsleep, 
         m17_inst_shutoff, m17_inst_mce, m17_inst_stbyp, m17_inst_wa_disable, 
         m17_inst_isolation_control_in, m18_inst_wen, m18_inst_ren, 
         m18_inst_async_rst, m18_inst_fastsleep, m18_inst_deepsleep, 
         m18_inst_shutoff, m18_inst_mce, m18_inst_stbyp, m18_inst_wa_disable, 
         m18_inst_isolation_control_in, m19_inst_wen, m19_inst_ren, 
         m19_inst_async_rst, m19_inst_fastsleep, m19_inst_deepsleep, 
         m19_inst_shutoff, m19_inst_mce, m19_inst_stbyp, m19_inst_wa_disable, 
         m19_inst_isolation_control_in, m20_inst_wen, m20_inst_ren, 
         m20_inst_async_rst, m20_inst_fastsleep, m20_inst_deepsleep, 
         m20_inst_shutoff, m20_inst_mce, m20_inst_stbyp, m20_inst_wa_disable, 
         m20_inst_isolation_control_in, m21_inst_wen, m21_inst_ren, 
         m21_inst_async_rst, m21_inst_fastsleep, m21_inst_deepsleep, 
         m21_inst_shutoff, m21_inst_mce, m21_inst_stbyp, m21_inst_wa_disable, 
         m21_inst_isolation_control_in, m22_inst_wen, m22_inst_ren, 
         m22_inst_async_rst, m22_inst_fastsleep, m22_inst_deepsleep, 
         m22_inst_shutoff, m22_inst_mce, m22_inst_stbyp, m22_inst_wa_disable, 
         m22_inst_isolation_control_in, m23_inst_wen, m23_inst_ren, 
         m23_inst_async_rst, m23_inst_fastsleep, m23_inst_deepsleep, 
         m23_inst_shutoff, m23_inst_mce, m23_inst_stbyp, m23_inst_wa_disable, 
         m23_inst_isolation_control_in, m24_inst_wen, m24_inst_ren, 
         m24_inst_async_rst, m24_inst_fastsleep, m24_inst_deepsleep, 
         m24_inst_shutoff, m24_inst_mce, m24_inst_stbyp, m24_inst_wa_disable, 
         m24_inst_isolation_control_in, m25_inst_wen, m25_inst_ren, 
         m25_inst_async_rst, m25_inst_fastsleep, m25_inst_deepsleep, 
         m25_inst_shutoff, m25_inst_mce, m25_inst_stbyp, m25_inst_wa_disable, 
         m25_inst_isolation_control_in, m26_inst_wen, m26_inst_ren, 
         m26_inst_async_rst, m26_inst_fastsleep, m26_inst_deepsleep, 
         m26_inst_shutoff, m26_inst_mce, m26_inst_stbyp, m26_inst_wa_disable, 
         m26_inst_isolation_control_in, m27_inst_wen, m27_inst_ren, 
         m27_inst_async_rst, m27_inst_fastsleep, m27_inst_deepsleep, 
         m27_inst_shutoff, m27_inst_mce, m27_inst_stbyp, m27_inst_wa_disable, 
         m27_inst_isolation_control_in, m28_inst_wen, m28_inst_ren, 
         m28_inst_async_rst, m28_inst_fastsleep, m28_inst_deepsleep, 
         m28_inst_shutoff, m28_inst_mce, m28_inst_stbyp, m28_inst_wa_disable, 
         m28_inst_isolation_control_in, m29_inst_wen, m29_inst_ren, 
         m29_inst_async_rst, m29_inst_fastsleep, m29_inst_deepsleep, 
         m29_inst_shutoff, m29_inst_mce, m29_inst_stbyp, m29_inst_wa_disable, 
         m29_inst_isolation_control_in, m30_inst_wen, m30_inst_ren, 
         m30_inst_async_rst, m30_inst_fastsleep, m30_inst_deepsleep, 
         m30_inst_shutoff, m30_inst_mce, m30_inst_stbyp, m30_inst_wa_disable, 
         m30_inst_isolation_control_in, m31_inst_wen, m31_inst_ren, 
         m31_inst_async_rst, m31_inst_fastsleep, m31_inst_deepsleep, 
         m31_inst_shutoff, m31_inst_mce, m31_inst_stbyp, m31_inst_wa_disable, 
         m31_inst_isolation_control_in, m32_inst_wen, m32_inst_ren, 
         m32_inst_async_rst, m32_inst_fastsleep, m32_inst_deepsleep, 
         m32_inst_shutoff, m32_inst_mce, m32_inst_stbyp, m32_inst_wa_disable, 
         m32_inst_isolation_control_in, m33_inst_wen, m33_inst_ren, 
         m33_inst_async_rst, m33_inst_fastsleep, m33_inst_deepsleep, 
         m33_inst_shutoff, m33_inst_mce, m33_inst_stbyp, m33_inst_wa_disable, 
         m33_inst_isolation_control_in, m34_inst_wen, m34_inst_ren, 
         m34_inst_async_rst, m34_inst_fastsleep, m34_inst_deepsleep, 
         m34_inst_shutoff, m34_inst_mce, m34_inst_stbyp, m34_inst_wa_disable, 
         m34_inst_isolation_control_in, m35_inst_wen, m35_inst_ren, 
         m35_inst_async_rst, m35_inst_fastsleep, m35_inst_deepsleep, 
         m35_inst_shutoff, m35_inst_mce, m35_inst_stbyp, m35_inst_wa_disable, 
         m35_inst_isolation_control_in, m36_inst_wen, m36_inst_ren, 
         m36_inst_async_rst, m36_inst_fastsleep, m36_inst_deepsleep, 
         m36_inst_shutoff, m36_inst_mce, m36_inst_stbyp, m36_inst_wa_disable, 
         m36_inst_isolation_control_in, m37_inst_wen, m37_inst_ren, 
         m37_inst_async_rst, m37_inst_fastsleep, m37_inst_deepsleep, 
         m37_inst_shutoff, m37_inst_mce, m37_inst_stbyp, m37_inst_wa_disable, 
         m37_inst_isolation_control_in, m38_inst_wen, m38_inst_ren, 
         m38_inst_async_rst, m38_inst_fastsleep, m38_inst_deepsleep, 
         m38_inst_shutoff, m38_inst_mce, m38_inst_stbyp, m38_inst_wa_disable, 
         m38_inst_isolation_control_in, m39_inst_wen, m39_inst_ren, 
         m39_inst_async_rst, m39_inst_fastsleep, m39_inst_deepsleep, 
         m39_inst_shutoff, m39_inst_mce, m39_inst_stbyp, m39_inst_wa_disable, 
         m39_inst_isolation_control_in, m40_inst_wen, m40_inst_ren, 
         m40_inst_async_rst, m40_inst_fastsleep, m40_inst_deepsleep, 
         m40_inst_shutoff, m40_inst_mce, m40_inst_stbyp, m40_inst_wa_disable, 
         m40_inst_isolation_control_in, reset, ijtag_select, si, capture_en, 
         shift_en, update_en, tck, bisr_si, bisr_se, bisr_clock, bisr_clear;
  output [71:0] m33_inst_q, m34_inst_q, m35_inst_q, m36_inst_q;
  output [31:0] m37_inst_q, m38_inst_q, m39_inst_q, m40_inst_q;
  output [21:0] m1_inst_q, m2_inst_q, m3_inst_q, m4_inst_q, m5_inst_q, 
                m6_inst_q, m7_inst_q, m8_inst_q, m9_inst_q, m10_inst_q, 
                m11_inst_q, m12_inst_q, m13_inst_q, m14_inst_q, m15_inst_q, 
                m16_inst_q, m17_inst_q, m18_inst_q, m19_inst_q, m20_inst_q, 
                m21_inst_q, m22_inst_q, m23_inst_q, m24_inst_q, m25_inst_q, 
                m26_inst_q, m27_inst_q, m28_inst_q, m29_inst_q, m30_inst_q, 
                m31_inst_q, m32_inst_q;
  output BIST_ON, BIST_DONE, BIST_GO, MBISTPG_STABLE, 
         m1_inst_dpslp_or_shutoffout, m1_inst_shutoffout, 
         m2_inst_dpslp_or_shutoffout, m2_inst_shutoffout, 
         m3_inst_dpslp_or_shutoffout, m3_inst_shutoffout, 
         m4_inst_dpslp_or_shutoffout, m4_inst_shutoffout, 
         m5_inst_dpslp_or_shutoffout, m5_inst_shutoffout, 
         m6_inst_dpslp_or_shutoffout, m6_inst_shutoffout, 
         m7_inst_dpslp_or_shutoffout, m7_inst_shutoffout, 
         m8_inst_dpslp_or_shutoffout, m8_inst_shutoffout, 
         m9_inst_dpslp_or_shutoffout, m9_inst_shutoffout, 
         m10_inst_dpslp_or_shutoffout, m10_inst_shutoffout, 
         m11_inst_dpslp_or_shutoffout, m11_inst_shutoffout, 
         m12_inst_dpslp_or_shutoffout, m12_inst_shutoffout, 
         m13_inst_dpslp_or_shutoffout, m13_inst_shutoffout, 
         m14_inst_dpslp_or_shutoffout, m14_inst_shutoffout, 
         m15_inst_dpslp_or_shutoffout, m15_inst_shutoffout, 
         m16_inst_dpslp_or_shutoffout, m16_inst_shutoffout, 
         m17_inst_dpslp_or_shutoffout, m17_inst_shutoffout, 
         m18_inst_dpslp_or_shutoffout, m18_inst_shutoffout, 
         m19_inst_dpslp_or_shutoffout, m19_inst_shutoffout, 
         m20_inst_dpslp_or_shutoffout, m20_inst_shutoffout, 
         m21_inst_dpslp_or_shutoffout, m21_inst_shutoffout, 
         m22_inst_dpslp_or_shutoffout, m22_inst_shutoffout, 
         m23_inst_dpslp_or_shutoffout, m23_inst_shutoffout, 
         m24_inst_dpslp_or_shutoffout, m24_inst_shutoffout, 
         m25_inst_dpslp_or_shutoffout, m25_inst_shutoffout, 
         m26_inst_dpslp_or_shutoffout, m26_inst_shutoffout, 
         m27_inst_dpslp_or_shutoffout, m27_inst_shutoffout, 
         m28_inst_dpslp_or_shutoffout, m28_inst_shutoffout, 
         m29_inst_dpslp_or_shutoffout, m29_inst_shutoffout, 
         m30_inst_dpslp_or_shutoffout, m30_inst_shutoffout, 
         m31_inst_dpslp_or_shutoffout, m31_inst_shutoffout, 
         m32_inst_dpslp_or_shutoffout, m32_inst_shutoffout, 
         m33_inst_dpslp_or_shutoffout, m33_inst_shutoffout, 
         m34_inst_dpslp_or_shutoffout, m34_inst_shutoffout, 
         m35_inst_dpslp_or_shutoffout, m35_inst_shutoffout, 
         m36_inst_dpslp_or_shutoffout, m36_inst_shutoffout, 
         m37_inst_dpslp_or_shutoffout, m37_inst_shutoffout, 
         m38_inst_dpslp_or_shutoffout, m38_inst_shutoffout, 
         m39_inst_dpslp_or_shutoffout, m39_inst_shutoffout, 
         m40_inst_dpslp_or_shutoffout, m40_inst_shutoffout, so, bisr_so;

  wire [71:0] din_ts25, din_ts26, din_ts27, din_ts28, m33_inst_q_ts1, 
              m34_inst_q_ts1, m35_inst_q_ts1, m36_inst_q_ts1;
  wire [31:0] din_ts29, din_ts30, din_ts31, din_ts33, m37_inst_q_ts1, 
              m38_inst_q_ts1, m39_inst_q_ts1, m40_inst_q_ts1;
  wire [25:0] c1_gate1_m33_bisr_inst_Q, c1_gate1_m34_bisr_inst_Q, 
              c1_gate1_m35_bisr_inst_Q, c1_gate1_m36_bisr_inst_Q;
  wire [21:0] din, din_ts1, din_ts2, din_ts3, din_ts4, din_ts5, din_ts6, 
              din_ts7, din_ts8, din_ts9, din_ts10, din_ts11, din_ts12, 
              din_ts13, din_ts14, din_ts15, din_ts16, din_ts17, din_ts18, 
              din_ts19, din_ts20, din_ts21, din_ts22, din_ts23, din_ts24, 
              din_ts32, din_ts34, din_ts35, din_ts36, din_ts37, din_ts38, 
              din_ts39, m10_inst_q_ts1, m11_inst_q_ts1, m12_inst_q_ts1, 
              m13_inst_q_ts1, m14_inst_q_ts1, m15_inst_q_ts1, m16_inst_q_ts1, 
              m17_inst_q_ts1, m18_inst_q_ts1, m19_inst_q_ts1, m1_inst_q_ts1, 
              m20_inst_q_ts1, m21_inst_q_ts1, m22_inst_q_ts1, m23_inst_q_ts1, 
              m24_inst_q_ts1, m25_inst_q_ts1, m26_inst_q_ts1, m27_inst_q_ts1, 
              m28_inst_q_ts1, m29_inst_q_ts1, m2_inst_q_ts1, m30_inst_q_ts1, 
              m31_inst_q_ts1, m32_inst_q_ts1, m3_inst_q_ts1, m4_inst_q_ts1, 
              m5_inst_q_ts1, m6_inst_q_ts1, m7_inst_q_ts1, m8_inst_q_ts1, 
              m9_inst_q_ts1, c1_gate1_m10_bisr_inst_Q, 
              c1_gate1_m11_bisr_inst_Q, c1_gate1_m12_bisr_inst_Q, 
              c1_gate1_m13_bisr_inst_Q, c1_gate1_m14_bisr_inst_Q, 
              c1_gate1_m15_bisr_inst_Q, c1_gate1_m16_bisr_inst_Q, 
              c1_gate1_m17_bisr_inst_Q, c1_gate1_m18_bisr_inst_Q, 
              c1_gate1_m19_bisr_inst_Q, c1_gate1_m1_bisr_inst_Q, 
              c1_gate1_m20_bisr_inst_Q, c1_gate1_m21_bisr_inst_Q, 
              c1_gate1_m22_bisr_inst_Q, c1_gate1_m23_bisr_inst_Q, 
              c1_gate1_m24_bisr_inst_Q, c1_gate1_m25_bisr_inst_Q, 
              c1_gate1_m26_bisr_inst_Q, c1_gate1_m27_bisr_inst_Q, 
              c1_gate1_m28_bisr_inst_Q, c1_gate1_m29_bisr_inst_Q, 
              c1_gate1_m2_bisr_inst_Q, c1_gate1_m30_bisr_inst_Q, 
              c1_gate1_m31_bisr_inst_Q, c1_gate1_m32_bisr_inst_Q, 
              c1_gate1_m37_bisr_inst_Q, c1_gate1_m38_bisr_inst_Q, 
              c1_gate1_m39_bisr_inst_Q, c1_gate1_m3_bisr_inst_Q, 
              c1_gate1_m40_bisr_inst_Q, c1_gate1_m4_bisr_inst_Q, 
              c1_gate1_m5_bisr_inst_Q, c1_gate1_m6_bisr_inst_Q, 
              c1_gate1_m7_bisr_inst_Q, c1_gate1_m8_bisr_inst_Q, 
              c1_gate1_m9_bisr_inst_Q;
  wire [9:0] adr, adr_ts1, adr_ts2, adr_ts3, adr_ts4, adr_ts5, adr_ts6, 
             adr_ts7, adr_ts8, adr_ts9, adr_ts10, adr_ts11, adr_ts12, adr_ts13, 
             adr_ts14, adr_ts15, adr_ts16, adr_ts17, adr_ts18, adr_ts19, 
             adr_ts20, adr_ts21, adr_ts22, adr_ts23, adr_ts24, adr_ts25, 
             adr_ts26, adr_ts27, adr_ts28, adr_ts32, adr_ts34, adr_ts35, 
             adr_ts36, adr_ts37, adr_ts38, adr_ts39;
  wire [8:0] adr_ts29, adr_ts30, adr_ts31, adr_ts33;
  wire [7:0] ALL_SROW0_FUSE_ADD_REG_ts25, ALL_SROW1_FUSE_ADD_REG_ts25, 
             ALL_SROW0_FUSE_ADD_REG_ts26, ALL_SROW1_FUSE_ADD_REG_ts26, 
             ALL_SROW0_FUSE_ADD_REG_ts27, ALL_SROW1_FUSE_ADD_REG_ts27, 
             ALL_SROW0_FUSE_ADD_REG_ts28, ALL_SROW1_FUSE_ADD_REG_ts28;
  wire [6:0] ALL_SROW0_FUSE_ADD_REG, ALL_SROW1_FUSE_ADD_REG, 
             ALL_SROW0_FUSE_ADD_REG_ts1, ALL_SROW1_FUSE_ADD_REG_ts1, 
             ALL_SROW0_FUSE_ADD_REG_ts2, ALL_SROW1_FUSE_ADD_REG_ts2, 
             ALL_SROW0_FUSE_ADD_REG_ts3, ALL_SROW1_FUSE_ADD_REG_ts3, 
             ALL_SROW0_FUSE_ADD_REG_ts4, ALL_SROW1_FUSE_ADD_REG_ts4, 
             ALL_SROW0_FUSE_ADD_REG_ts5, ALL_SROW1_FUSE_ADD_REG_ts5, 
             ALL_SROW0_FUSE_ADD_REG_ts6, ALL_SROW1_FUSE_ADD_REG_ts6, 
             ALL_SROW0_FUSE_ADD_REG_ts7, ALL_SROW1_FUSE_ADD_REG_ts7, 
             ALL_SROW0_FUSE_ADD_REG_ts8, ALL_SROW1_FUSE_ADD_REG_ts8, 
             ALL_SROW0_FUSE_ADD_REG_ts9, ALL_SROW1_FUSE_ADD_REG_ts9, 
             ALL_SROW0_FUSE_ADD_REG_ts10, ALL_SROW1_FUSE_ADD_REG_ts10, 
             ALL_SROW0_FUSE_ADD_REG_ts11, ALL_SROW1_FUSE_ADD_REG_ts11, 
             ALL_SROW0_FUSE_ADD_REG_ts12, ALL_SROW1_FUSE_ADD_REG_ts12, 
             ALL_SROW0_FUSE_ADD_REG_ts13, ALL_SROW1_FUSE_ADD_REG_ts13, 
             ALL_SROW0_FUSE_ADD_REG_ts14, ALL_SROW1_FUSE_ADD_REG_ts14, 
             ALL_SROW0_FUSE_ADD_REG_ts15, ALL_SROW1_FUSE_ADD_REG_ts15, 
             ALL_SROW0_FUSE_ADD_REG_ts16, ALL_SROW1_FUSE_ADD_REG_ts16, 
             ALL_SROW0_FUSE_ADD_REG_ts17, ALL_SROW1_FUSE_ADD_REG_ts17, 
             ALL_SROW0_FUSE_ADD_REG_ts18, ALL_SROW1_FUSE_ADD_REG_ts18, 
             ALL_SROW0_FUSE_ADD_REG_ts19, ALL_SROW1_FUSE_ADD_REG_ts19, 
             ALL_SROW0_FUSE_ADD_REG_ts20, ALL_SROW1_FUSE_ADD_REG_ts20, 
             ALL_SROW0_FUSE_ADD_REG_ts21, ALL_SROW1_FUSE_ADD_REG_ts21, 
             ALL_SROW0_FUSE_ADD_REG_ts22, ALL_SROW1_FUSE_ADD_REG_ts22, 
             ALL_SROW0_FUSE_ADD_REG_ts23, ALL_SROW1_FUSE_ADD_REG_ts23, 
             ALL_SROW0_FUSE_ADD_REG_ts24, ALL_SROW1_FUSE_ADD_REG_ts24, 
             All_SCOL0_FUSE_REG_ts25, All_SCOL0_FUSE_REG_ts26, 
             All_SCOL0_FUSE_REG_ts27, All_SCOL0_FUSE_REG_ts28, 
             ALL_SROW0_FUSE_ADD_REG_ts29, ALL_SROW1_FUSE_ADD_REG_ts29, 
             ALL_SROW0_FUSE_ADD_REG_ts30, ALL_SROW1_FUSE_ADD_REG_ts30, 
             ALL_SROW0_FUSE_ADD_REG_ts31, ALL_SROW1_FUSE_ADD_REG_ts31, 
             ALL_SROW0_FUSE_ADD_REG_ts32, ALL_SROW1_FUSE_ADD_REG_ts32, 
             ALL_SROW0_FUSE_ADD_REG_ts33, ALL_SROW1_FUSE_ADD_REG_ts33, 
             ALL_SROW0_FUSE_ADD_REG_ts34, ALL_SROW1_FUSE_ADD_REG_ts34, 
             ALL_SROW0_FUSE_ADD_REG_ts35, ALL_SROW1_FUSE_ADD_REG_ts35, 
             ALL_SROW0_FUSE_ADD_REG_ts36, ALL_SROW1_FUSE_ADD_REG_ts36, 
             ALL_SROW0_FUSE_ADD_REG_ts37, ALL_SROW1_FUSE_ADD_REG_ts37, 
             ALL_SROW0_FUSE_ADD_REG_ts38, ALL_SROW1_FUSE_ADD_REG_ts38, 
             ALL_SROW0_FUSE_ADD_REG_ts39, ALL_SROW1_FUSE_ADD_REG_ts39;
  wire [4:0] All_SCOL0_FUSE_REG, All_SCOL0_FUSE_REG_ts1, 
             All_SCOL0_FUSE_REG_ts2, All_SCOL0_FUSE_REG_ts3, 
             All_SCOL0_FUSE_REG_ts4, All_SCOL0_FUSE_REG_ts5, 
             All_SCOL0_FUSE_REG_ts6, All_SCOL0_FUSE_REG_ts7, 
             All_SCOL0_FUSE_REG_ts8, All_SCOL0_FUSE_REG_ts9, 
             All_SCOL0_FUSE_REG_ts10, All_SCOL0_FUSE_REG_ts11, 
             All_SCOL0_FUSE_REG_ts12, All_SCOL0_FUSE_REG_ts13, 
             All_SCOL0_FUSE_REG_ts14, All_SCOL0_FUSE_REG_ts15, 
             All_SCOL0_FUSE_REG_ts16, All_SCOL0_FUSE_REG_ts17, 
             All_SCOL0_FUSE_REG_ts18, All_SCOL0_FUSE_REG_ts19, 
             All_SCOL0_FUSE_REG_ts20, All_SCOL0_FUSE_REG_ts21, 
             All_SCOL0_FUSE_REG_ts22, All_SCOL0_FUSE_REG_ts23, 
             All_SCOL0_FUSE_REG_ts24, All_SCOL0_FUSE_REG_ts29, 
             All_SCOL0_FUSE_REG_ts30, All_SCOL0_FUSE_REG_ts31, 
             All_SCOL0_FUSE_REG_ts32, All_SCOL0_FUSE_REG_ts33, 
             All_SCOL0_FUSE_REG_ts34, All_SCOL0_FUSE_REG_ts35, 
             All_SCOL0_FUSE_REG_ts36, All_SCOL0_FUSE_REG_ts37, 
             All_SCOL0_FUSE_REG_ts38, All_SCOL0_FUSE_REG_ts39;
  wire [0:0] toBist, bistEn;
  wire BIRA_EN, PRESERVE_FUSE_REGISTER, CHECK_REPAIR_NEEDED, BIST_HOLD, 
       BIST_SETUP, BIST_SETUP_ts1, BIST_SETUP_ts2, BIST_SELECT_TEST_DATA, 
       to_controllers_tck, mcp_bounding_to_en, scan_to_en, memory_bypass_to_en, 
       ltest_to_en, BIST_ALGO_MODE0, BIST_ALGO_MODE1, ENABLE_MEM_RESET, 
       REDUCED_ADDRESS_COUNT, MEM_ARRAY_DUMP_MODE, BIST_DIAG_EN, 
       BIST_CLEAR_BIRA, BIST_COLLAR_DIAG_EN, BIST_COLLAR_BIRA_EN, 
       PriorityColumn, BIST_SHIFT_BIRA_COLLAR, BIST_ASYNC_RESET, 
       MEM0_BIST_COLLAR_SI, MEM1_BIST_COLLAR_SI, MEM2_BIST_COLLAR_SI, 
       MEM3_BIST_COLLAR_SI, MEM4_BIST_COLLAR_SI, MEM5_BIST_COLLAR_SI, 
       MEM6_BIST_COLLAR_SI, MEM7_BIST_COLLAR_SI, MEM8_BIST_COLLAR_SI, 
       MEM9_BIST_COLLAR_SI, MEM10_BIST_COLLAR_SI, MEM11_BIST_COLLAR_SI, 
       MEM12_BIST_COLLAR_SI, MEM13_BIST_COLLAR_SI, MEM14_BIST_COLLAR_SI, 
       MEM15_BIST_COLLAR_SI, MEM16_BIST_COLLAR_SI, MEM17_BIST_COLLAR_SI, 
       MEM18_BIST_COLLAR_SI, MEM19_BIST_COLLAR_SI, MEM20_BIST_COLLAR_SI, 
       MEM21_BIST_COLLAR_SI, MEM22_BIST_COLLAR_SI, MEM23_BIST_COLLAR_SI, 
       MEM24_BIST_COLLAR_SI, MEM25_BIST_COLLAR_SI, MEM26_BIST_COLLAR_SI, 
       MEM27_BIST_COLLAR_SI, MEM28_BIST_COLLAR_SI, MEM29_BIST_COLLAR_SI, 
       MEM30_BIST_COLLAR_SI, MEM31_BIST_COLLAR_SI, MEM32_BIST_COLLAR_SI, 
       MEM33_BIST_COLLAR_SI, MEM34_BIST_COLLAR_SI, MEM35_BIST_COLLAR_SI, 
       MEM36_BIST_COLLAR_SI, MEM37_BIST_COLLAR_SI, MEM38_BIST_COLLAR_SI, 
       MEM39_BIST_COLLAR_SI, MBISTPG_SO, BIST_SO, BIST_SO_ts1, BIST_SO_ts2, 
       BIST_SO_ts3, BIST_SO_ts4, BIST_SO_ts5, BIST_SO_ts6, BIST_SO_ts7, 
       BIST_SO_ts8, BIST_SO_ts9, BIST_SO_ts10, BIST_SO_ts11, BIST_SO_ts12, 
       BIST_SO_ts13, BIST_SO_ts14, BIST_SO_ts15, BIST_SO_ts16, BIST_SO_ts17, 
       BIST_SO_ts18, BIST_SO_ts19, BIST_SO_ts20, BIST_SO_ts21, BIST_SO_ts22, 
       BIST_SO_ts23, BIST_SO_ts24, BIST_SO_ts25, BIST_SO_ts26, BIST_SO_ts27, 
       BIST_SO_ts28, BIST_SO_ts29, BIST_SO_ts30, BIST_SO_ts31, BIST_SO_ts32, 
       BIST_SO_ts33, BIST_SO_ts34, BIST_SO_ts35, BIST_SO_ts36, BIST_SO_ts37, 
       BIST_SO_ts38, BIST_SO_ts39, BIST_GO_ts1, BIST_GO_ts2, BIST_GO_ts3, 
       BIST_GO_ts4, BIST_GO_ts5, BIST_GO_ts6, BIST_GO_ts7, BIST_GO_ts8, 
       BIST_GO_ts9, BIST_GO_ts10, BIST_GO_ts11, BIST_GO_ts12, BIST_GO_ts13, 
       BIST_GO_ts14, BIST_GO_ts15, BIST_GO_ts16, BIST_GO_ts17, BIST_GO_ts18, 
       BIST_GO_ts19, BIST_GO_ts20, BIST_GO_ts21, BIST_GO_ts22, BIST_GO_ts23, 
       BIST_GO_ts24, BIST_GO_ts25, BIST_GO_ts26, BIST_GO_ts27, BIST_GO_ts28, 
       BIST_GO_ts29, BIST_GO_ts30, BIST_GO_ts31, BIST_GO_ts32, BIST_GO_ts33, 
       BIST_GO_ts34, BIST_GO_ts35, BIST_GO_ts36, BIST_GO_ts37, BIST_GO_ts38, 
       BIST_GO_ts39, BIST_GO_ts40, FL_CNT_MODE0, FL_CNT_MODE1, 
       BIST_WRITEENABLE, BIST_READENABLE, BIST_CMP, INCLUDE_MEM_RESULTS_REG, 
       BIST_COL_ADD, BIST_COL_ADD_ts1, BIST_COL_ADD_ts2, BIST_ROW_ADD, 
       BIST_ROW_ADD_ts1, BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts4, 
       BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts7, BIST_COLLAR_EN0, 
       BIST_COLLAR_EN1, BIST_COLLAR_EN2, BIST_COLLAR_EN3, BIST_COLLAR_EN4, 
       BIST_COLLAR_EN5, BIST_COLLAR_EN6, BIST_COLLAR_EN7, BIST_COLLAR_EN8, 
       BIST_COLLAR_EN9, BIST_COLLAR_EN10, BIST_COLLAR_EN11, BIST_COLLAR_EN12, 
       BIST_COLLAR_EN13, BIST_COLLAR_EN14, BIST_COLLAR_EN15, BIST_COLLAR_EN16, 
       BIST_COLLAR_EN17, BIST_COLLAR_EN18, BIST_COLLAR_EN19, BIST_COLLAR_EN20, 
       BIST_COLLAR_EN21, BIST_COLLAR_EN22, BIST_COLLAR_EN23, BIST_COLLAR_EN24, 
       BIST_COLLAR_EN25, BIST_COLLAR_EN26, BIST_COLLAR_EN27, BIST_COLLAR_EN28, 
       BIST_COLLAR_EN29, BIST_COLLAR_EN30, BIST_COLLAR_EN31, BIST_COLLAR_EN32, 
       BIST_COLLAR_EN33, BIST_COLLAR_EN34, BIST_COLLAR_EN35, BIST_COLLAR_EN36, 
       BIST_COLLAR_EN37, BIST_COLLAR_EN38, BIST_COLLAR_EN39, 
       BIST_RUN_TO_COLLAR0, BIST_RUN_TO_COLLAR1, BIST_RUN_TO_COLLAR2, 
       BIST_RUN_TO_COLLAR3, BIST_RUN_TO_COLLAR4, BIST_RUN_TO_COLLAR5, 
       BIST_RUN_TO_COLLAR6, BIST_RUN_TO_COLLAR7, BIST_RUN_TO_COLLAR8, 
       BIST_RUN_TO_COLLAR9, BIST_RUN_TO_COLLAR10, BIST_RUN_TO_COLLAR11, 
       BIST_RUN_TO_COLLAR12, BIST_RUN_TO_COLLAR13, BIST_RUN_TO_COLLAR14, 
       BIST_RUN_TO_COLLAR15, BIST_RUN_TO_COLLAR16, BIST_RUN_TO_COLLAR17, 
       BIST_RUN_TO_COLLAR18, BIST_RUN_TO_COLLAR19, BIST_RUN_TO_COLLAR20, 
       BIST_RUN_TO_COLLAR21, BIST_RUN_TO_COLLAR22, BIST_RUN_TO_COLLAR23, 
       BIST_RUN_TO_COLLAR24, BIST_RUN_TO_COLLAR25, BIST_RUN_TO_COLLAR26, 
       BIST_RUN_TO_COLLAR27, BIST_RUN_TO_COLLAR28, BIST_RUN_TO_COLLAR29, 
       BIST_RUN_TO_COLLAR30, BIST_RUN_TO_COLLAR31, BIST_RUN_TO_COLLAR32, 
       BIST_RUN_TO_COLLAR33, BIST_RUN_TO_COLLAR34, BIST_RUN_TO_COLLAR35, 
       BIST_RUN_TO_COLLAR36, BIST_RUN_TO_COLLAR37, BIST_RUN_TO_COLLAR38, 
       BIST_RUN_TO_COLLAR39, to_interfaces_tck, BIST_TESTDATA_SELECT_TO_COLLAR, 
       BIST_WRITE_DATA, BIST_WRITE_DATA_ts1, BIST_WRITE_DATA_ts2, 
       BIST_WRITE_DATA_ts3, BIST_EXPECT_DATA, BIST_EXPECT_DATA_ts1, 
       BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts3, CHKBCI_PHASE, 
       BIST_SHIFT_COLLAR, BIST_COLLAR_SETUP, BIST_CLEAR_DEFAULT, BIST_CLEAR, 
       BIST_COLLAR_OPSET_SELECT, BIST_COLLAR_HOLD, FREEZE_STOP_ERROR, 
       ERROR_CNT_ZERO, MBISTPG_RESET_REG_SETUP2, wen, wen_ts1, wen_ts2, 
       wen_ts3, wen_ts4, wen_ts5, wen_ts6, wen_ts7, wen_ts8, wen_ts9, wen_ts10, 
       wen_ts11, wen_ts12, wen_ts13, wen_ts14, wen_ts15, wen_ts16, wen_ts17, 
       wen_ts18, wen_ts19, wen_ts20, wen_ts21, wen_ts22, wen_ts23, wen_ts24, 
       wen_ts25, wen_ts26, wen_ts27, wen_ts28, wen_ts29, wen_ts30, wen_ts31, 
       wen_ts32, wen_ts33, wen_ts34, wen_ts35, wen_ts36, wen_ts37, wen_ts38, 
       wen_ts39, ren, ren_ts1, ren_ts2, ren_ts3, ren_ts4, ren_ts5, ren_ts6, 
       ren_ts7, ren_ts8, ren_ts9, ren_ts10, ren_ts11, ren_ts12, ren_ts13, 
       ren_ts14, ren_ts15, ren_ts16, ren_ts17, ren_ts18, ren_ts19, ren_ts20, 
       ren_ts21, ren_ts22, ren_ts23, ren_ts24, ren_ts25, ren_ts26, ren_ts27, 
       ren_ts28, ren_ts29, ren_ts30, ren_ts31, ren_ts32, ren_ts33, ren_ts34, 
       ren_ts35, ren_ts36, ren_ts37, ren_ts38, ren_ts39, bisr_so_ts1, 
       c1_gate1_m10_bisr_inst_SO, c1_gate1_m11_bisr_inst_SO, 
       c1_gate1_m12_bisr_inst_SO, c1_gate1_m13_bisr_inst_SO, 
       c1_gate1_m14_bisr_inst_SO, c1_gate1_m15_bisr_inst_SO, 
       c1_gate1_m16_bisr_inst_SO, c1_gate1_m17_bisr_inst_SO, 
       c1_gate1_m18_bisr_inst_SO, c1_gate1_m19_bisr_inst_SO, 
       c1_gate1_m1_bisr_inst_SO, c1_gate1_m20_bisr_inst_SO, 
       c1_gate1_m21_bisr_inst_SO, c1_gate1_m22_bisr_inst_SO, 
       c1_gate1_m23_bisr_inst_SO, c1_gate1_m24_bisr_inst_SO, 
       c1_gate1_m25_bisr_inst_SO, c1_gate1_m26_bisr_inst_SO, 
       c1_gate1_m27_bisr_inst_SO, c1_gate1_m28_bisr_inst_SO, 
       c1_gate1_m29_bisr_inst_SO, c1_gate1_m2_bisr_inst_SO, 
       c1_gate1_m30_bisr_inst_SO, c1_gate1_m31_bisr_inst_SO, 
       c1_gate1_m32_bisr_inst_SO, c1_gate1_m33_bisr_inst_SO, 
       c1_gate1_m34_bisr_inst_SO, c1_gate1_m35_bisr_inst_SO, 
       c1_gate1_m36_bisr_inst_SO, c1_gate1_m37_bisr_inst_SO, 
       c1_gate1_m38_bisr_inst_SO, c1_gate1_m39_bisr_inst_SO, 
       c1_gate1_m3_bisr_inst_SO, c1_gate1_m4_bisr_inst_SO, 
       c1_gate1_m5_bisr_inst_SO, c1_gate1_m6_bisr_inst_SO, 
       c1_gate1_m7_bisr_inst_SO, c1_gate1_m8_bisr_inst_SO, 
       c1_gate1_m9_bisr_inst_SO, ALL_SROW0_ALLOC_REG, ALL_SROW1_ALLOC_REG, 
       All_SCOL0_ALLOC_REG, ALL_SROW0_ALLOC_REG_ts1, ALL_SROW1_ALLOC_REG_ts1, 
       All_SCOL0_ALLOC_REG_ts1, ALL_SROW0_ALLOC_REG_ts2, 
       ALL_SROW1_ALLOC_REG_ts2, All_SCOL0_ALLOC_REG_ts2, 
       ALL_SROW0_ALLOC_REG_ts3, ALL_SROW1_ALLOC_REG_ts3, 
       All_SCOL0_ALLOC_REG_ts3, ALL_SROW0_ALLOC_REG_ts4, 
       ALL_SROW1_ALLOC_REG_ts4, All_SCOL0_ALLOC_REG_ts4, 
       ALL_SROW0_ALLOC_REG_ts5, ALL_SROW1_ALLOC_REG_ts5, 
       All_SCOL0_ALLOC_REG_ts5, ALL_SROW0_ALLOC_REG_ts6, 
       ALL_SROW1_ALLOC_REG_ts6, All_SCOL0_ALLOC_REG_ts6, 
       ALL_SROW0_ALLOC_REG_ts7, ALL_SROW1_ALLOC_REG_ts7, 
       All_SCOL0_ALLOC_REG_ts7, ALL_SROW0_ALLOC_REG_ts8, 
       ALL_SROW1_ALLOC_REG_ts8, All_SCOL0_ALLOC_REG_ts8, 
       ALL_SROW0_ALLOC_REG_ts9, ALL_SROW1_ALLOC_REG_ts9, 
       All_SCOL0_ALLOC_REG_ts9, ALL_SROW0_ALLOC_REG_ts10, 
       ALL_SROW1_ALLOC_REG_ts10, All_SCOL0_ALLOC_REG_ts10, 
       ALL_SROW0_ALLOC_REG_ts11, ALL_SROW1_ALLOC_REG_ts11, 
       All_SCOL0_ALLOC_REG_ts11, ALL_SROW0_ALLOC_REG_ts12, 
       ALL_SROW1_ALLOC_REG_ts12, All_SCOL0_ALLOC_REG_ts12, 
       ALL_SROW0_ALLOC_REG_ts13, ALL_SROW1_ALLOC_REG_ts13, 
       All_SCOL0_ALLOC_REG_ts13, ALL_SROW0_ALLOC_REG_ts14, 
       ALL_SROW1_ALLOC_REG_ts14, All_SCOL0_ALLOC_REG_ts14, 
       ALL_SROW0_ALLOC_REG_ts15, ALL_SROW1_ALLOC_REG_ts15, 
       All_SCOL0_ALLOC_REG_ts15, ALL_SROW0_ALLOC_REG_ts16, 
       ALL_SROW1_ALLOC_REG_ts16, All_SCOL0_ALLOC_REG_ts16, 
       ALL_SROW0_ALLOC_REG_ts17, ALL_SROW1_ALLOC_REG_ts17, 
       All_SCOL0_ALLOC_REG_ts17, ALL_SROW0_ALLOC_REG_ts18, 
       ALL_SROW1_ALLOC_REG_ts18, All_SCOL0_ALLOC_REG_ts18, 
       ALL_SROW0_ALLOC_REG_ts19, ALL_SROW1_ALLOC_REG_ts19, 
       All_SCOL0_ALLOC_REG_ts19, ALL_SROW0_ALLOC_REG_ts20, 
       ALL_SROW1_ALLOC_REG_ts20, All_SCOL0_ALLOC_REG_ts20, 
       ALL_SROW0_ALLOC_REG_ts21, ALL_SROW1_ALLOC_REG_ts21, 
       All_SCOL0_ALLOC_REG_ts21, ALL_SROW0_ALLOC_REG_ts22, 
       ALL_SROW1_ALLOC_REG_ts22, All_SCOL0_ALLOC_REG_ts22, 
       ALL_SROW0_ALLOC_REG_ts23, ALL_SROW1_ALLOC_REG_ts23, 
       All_SCOL0_ALLOC_REG_ts23, ALL_SROW0_ALLOC_REG_ts24, 
       ALL_SROW1_ALLOC_REG_ts24, All_SCOL0_ALLOC_REG_ts24, 
       ALL_SROW0_ALLOC_REG_ts25, ALL_SROW1_ALLOC_REG_ts25, 
       All_SCOL0_ALLOC_REG_ts25, ALL_SROW0_ALLOC_REG_ts26, 
       ALL_SROW1_ALLOC_REG_ts26, All_SCOL0_ALLOC_REG_ts26, 
       ALL_SROW0_ALLOC_REG_ts27, ALL_SROW1_ALLOC_REG_ts27, 
       All_SCOL0_ALLOC_REG_ts27, ALL_SROW0_ALLOC_REG_ts28, 
       ALL_SROW1_ALLOC_REG_ts28, All_SCOL0_ALLOC_REG_ts28, 
       ALL_SROW0_ALLOC_REG_ts29, ALL_SROW1_ALLOC_REG_ts29, 
       All_SCOL0_ALLOC_REG_ts29, ALL_SROW0_ALLOC_REG_ts30, 
       ALL_SROW1_ALLOC_REG_ts30, All_SCOL0_ALLOC_REG_ts30, 
       ALL_SROW0_ALLOC_REG_ts31, ALL_SROW1_ALLOC_REG_ts31, 
       All_SCOL0_ALLOC_REG_ts31, ALL_SROW0_ALLOC_REG_ts32, 
       ALL_SROW1_ALLOC_REG_ts32, All_SCOL0_ALLOC_REG_ts32, 
       ALL_SROW0_ALLOC_REG_ts33, ALL_SROW1_ALLOC_REG_ts33, 
       All_SCOL0_ALLOC_REG_ts33, ALL_SROW0_ALLOC_REG_ts34, 
       ALL_SROW1_ALLOC_REG_ts34, All_SCOL0_ALLOC_REG_ts34, 
       ALL_SROW0_ALLOC_REG_ts35, ALL_SROW1_ALLOC_REG_ts35, 
       All_SCOL0_ALLOC_REG_ts35, ALL_SROW0_ALLOC_REG_ts36, 
       ALL_SROW1_ALLOC_REG_ts36, All_SCOL0_ALLOC_REG_ts36, 
       ALL_SROW0_ALLOC_REG_ts37, ALL_SROW1_ALLOC_REG_ts37, 
       All_SCOL0_ALLOC_REG_ts37, ALL_SROW0_ALLOC_REG_ts38, 
       ALL_SROW1_ALLOC_REG_ts38, All_SCOL0_ALLOC_REG_ts38, 
       ALL_SROW0_ALLOC_REG_ts39, ALL_SROW1_ALLOC_REG_ts39, 
       All_SCOL0_ALLOC_REG_ts39;

  assign bisr_so_ts1 = bisr_si;
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m1_inst(
      .row_repair_in({m1_inst_row_repair_in[25:21], 
      c1_gate1_m1_bisr_inst_Q[15:8], m1_inst_row_repair_in[12:8], 
      c1_gate1_m1_bisr_inst_Q[7:0]}), .col_repair_in({
      m1_inst_col_repair_in[12:6], c1_gate1_m1_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts10), .ren(ren_ts10), .async_rst(m1_inst_async_rst), .fastsleep(m1_inst_fastsleep), 
      .deepsleep(m1_inst_deepsleep), .sbc(m1_inst_sbc), .shutoff(m1_inst_shutoff), 
      .mce(m1_inst_mce), .stbyp(m1_inst_stbyp), .rmce(m1_inst_rmce), .wmce(m1_inst_wmce), 
      .wpulse(m1_inst_wpulse), .wa_disable(m1_inst_wa_disable), .wa(m1_inst_wa), 
      .ra(m1_inst_ra), .global_rrow_en_in(m1_inst_global_rrow_en_in), .isolation_control_in(m1_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m1_inst_dpslp_or_shutoffout), .shutoffout(m1_inst_shutoffout), 
      .adr(adr_ts10), .din(din_ts10), .q(m1_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m2_inst(
      .row_repair_in({m2_inst_row_repair_in[25:21], 
      c1_gate1_m2_bisr_inst_Q[15:8], m2_inst_row_repair_in[12:8], 
      c1_gate1_m2_bisr_inst_Q[7:0]}), .col_repair_in({
      m2_inst_col_repair_in[12:6], c1_gate1_m2_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts21), .ren(ren_ts21), .async_rst(m2_inst_async_rst), .fastsleep(m2_inst_fastsleep), 
      .deepsleep(m2_inst_deepsleep), .sbc(m2_inst_sbc), .shutoff(m2_inst_shutoff), 
      .mce(m2_inst_mce), .stbyp(m2_inst_stbyp), .rmce(m2_inst_rmce), .wmce(m2_inst_wmce), 
      .wpulse(m2_inst_wpulse), .wa_disable(m2_inst_wa_disable), .wa(m2_inst_wa), 
      .ra(m2_inst_ra), .global_rrow_en_in(m2_inst_global_rrow_en_in), .isolation_control_in(m2_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m2_inst_dpslp_or_shutoffout), .shutoffout(m2_inst_shutoffout), 
      .adr(adr_ts21), .din(din_ts21), .q(m2_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m3_inst(
      .row_repair_in({m3_inst_row_repair_in[25:21], 
      c1_gate1_m3_bisr_inst_Q[15:8], m3_inst_row_repair_in[12:8], 
      c1_gate1_m3_bisr_inst_Q[7:0]}), .col_repair_in({
      m3_inst_col_repair_in[12:6], c1_gate1_m3_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts32), .ren(ren_ts32), .async_rst(m3_inst_async_rst), .fastsleep(m3_inst_fastsleep), 
      .deepsleep(m3_inst_deepsleep), .sbc(m3_inst_sbc), .shutoff(m3_inst_shutoff), 
      .mce(m3_inst_mce), .stbyp(m3_inst_stbyp), .rmce(m3_inst_rmce), .wmce(m3_inst_wmce), 
      .wpulse(m3_inst_wpulse), .wa_disable(m3_inst_wa_disable), .wa(m3_inst_wa), 
      .ra(m3_inst_ra), .global_rrow_en_in(m3_inst_global_rrow_en_in), .isolation_control_in(m3_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m3_inst_dpslp_or_shutoffout), .shutoffout(m3_inst_shutoffout), 
      .adr(adr_ts32), .din(din_ts32), .q(m3_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m4_inst(
      .row_repair_in({m4_inst_row_repair_in[25:21], 
      c1_gate1_m4_bisr_inst_Q[15:8], m4_inst_row_repair_in[12:8], 
      c1_gate1_m4_bisr_inst_Q[7:0]}), .col_repair_in({
      m4_inst_col_repair_in[12:6], c1_gate1_m4_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts34), .ren(ren_ts34), .async_rst(m4_inst_async_rst), .fastsleep(m4_inst_fastsleep), 
      .deepsleep(m4_inst_deepsleep), .sbc(m4_inst_sbc), .shutoff(m4_inst_shutoff), 
      .mce(m4_inst_mce), .stbyp(m4_inst_stbyp), .rmce(m4_inst_rmce), .wmce(m4_inst_wmce), 
      .wpulse(m4_inst_wpulse), .wa_disable(m4_inst_wa_disable), .wa(m4_inst_wa), 
      .ra(m4_inst_ra), .global_rrow_en_in(m4_inst_global_rrow_en_in), .isolation_control_in(m4_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m4_inst_dpslp_or_shutoffout), .shutoffout(m4_inst_shutoffout), 
      .adr(adr_ts34), .din(din_ts34), .q(m4_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m5_inst(
      .row_repair_in({m5_inst_row_repair_in[25:21], 
      c1_gate1_m5_bisr_inst_Q[15:8], m5_inst_row_repair_in[12:8], 
      c1_gate1_m5_bisr_inst_Q[7:0]}), .col_repair_in({
      m5_inst_col_repair_in[12:6], c1_gate1_m5_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts35), .ren(ren_ts35), .async_rst(m5_inst_async_rst), .fastsleep(m5_inst_fastsleep), 
      .deepsleep(m5_inst_deepsleep), .sbc(m5_inst_sbc), .shutoff(m5_inst_shutoff), 
      .mce(m5_inst_mce), .stbyp(m5_inst_stbyp), .rmce(m5_inst_rmce), .wmce(m5_inst_wmce), 
      .wpulse(m5_inst_wpulse), .wa_disable(m5_inst_wa_disable), .wa(m5_inst_wa), 
      .ra(m5_inst_ra), .global_rrow_en_in(m5_inst_global_rrow_en_in), .isolation_control_in(m5_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m5_inst_dpslp_or_shutoffout), .shutoffout(m5_inst_shutoffout), 
      .adr(adr_ts35), .din(din_ts35), .q(m5_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m6_inst(
      .row_repair_in({m6_inst_row_repair_in[25:21], 
      c1_gate1_m6_bisr_inst_Q[15:8], m6_inst_row_repair_in[12:8], 
      c1_gate1_m6_bisr_inst_Q[7:0]}), .col_repair_in({
      m6_inst_col_repair_in[12:6], c1_gate1_m6_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts36), .ren(ren_ts36), .async_rst(m6_inst_async_rst), .fastsleep(m6_inst_fastsleep), 
      .deepsleep(m6_inst_deepsleep), .sbc(m6_inst_sbc), .shutoff(m6_inst_shutoff), 
      .mce(m6_inst_mce), .stbyp(m6_inst_stbyp), .rmce(m6_inst_rmce), .wmce(m6_inst_wmce), 
      .wpulse(m6_inst_wpulse), .wa_disable(m6_inst_wa_disable), .wa(m6_inst_wa), 
      .ra(m6_inst_ra), .global_rrow_en_in(m6_inst_global_rrow_en_in), .isolation_control_in(m6_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m6_inst_dpslp_or_shutoffout), .shutoffout(m6_inst_shutoffout), 
      .adr(adr_ts36), .din(din_ts36), .q(m6_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m7_inst(
      .row_repair_in({m7_inst_row_repair_in[25:21], 
      c1_gate1_m7_bisr_inst_Q[15:8], m7_inst_row_repair_in[12:8], 
      c1_gate1_m7_bisr_inst_Q[7:0]}), .col_repair_in({
      m7_inst_col_repair_in[12:6], c1_gate1_m7_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts37), .ren(ren_ts37), .async_rst(m7_inst_async_rst), .fastsleep(m7_inst_fastsleep), 
      .deepsleep(m7_inst_deepsleep), .sbc(m7_inst_sbc), .shutoff(m7_inst_shutoff), 
      .mce(m7_inst_mce), .stbyp(m7_inst_stbyp), .rmce(m7_inst_rmce), .wmce(m7_inst_wmce), 
      .wpulse(m7_inst_wpulse), .wa_disable(m7_inst_wa_disable), .wa(m7_inst_wa), 
      .ra(m7_inst_ra), .global_rrow_en_in(m7_inst_global_rrow_en_in), .isolation_control_in(m7_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m7_inst_dpslp_or_shutoffout), .shutoffout(m7_inst_shutoffout), 
      .adr(adr_ts37), .din(din_ts37), .q(m7_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m8_inst(
      .row_repair_in({m8_inst_row_repair_in[25:21], 
      c1_gate1_m8_bisr_inst_Q[15:8], m8_inst_row_repair_in[12:8], 
      c1_gate1_m8_bisr_inst_Q[7:0]}), .col_repair_in({
      m8_inst_col_repair_in[12:6], c1_gate1_m8_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts38), .ren(ren_ts38), .async_rst(m8_inst_async_rst), .fastsleep(m8_inst_fastsleep), 
      .deepsleep(m8_inst_deepsleep), .sbc(m8_inst_sbc), .shutoff(m8_inst_shutoff), 
      .mce(m8_inst_mce), .stbyp(m8_inst_stbyp), .rmce(m8_inst_rmce), .wmce(m8_inst_wmce), 
      .wpulse(m8_inst_wpulse), .wa_disable(m8_inst_wa_disable), .wa(m8_inst_wa), 
      .ra(m8_inst_ra), .global_rrow_en_in(m8_inst_global_rrow_en_in), .isolation_control_in(m8_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m8_inst_dpslp_or_shutoffout), .shutoffout(m8_inst_shutoffout), 
      .adr(adr_ts38), .din(din_ts38), .q(m8_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m9_inst(
      .row_repair_in({m9_inst_row_repair_in[25:21], 
      c1_gate1_m9_bisr_inst_Q[15:8], m9_inst_row_repair_in[12:8], 
      c1_gate1_m9_bisr_inst_Q[7:0]}), .col_repair_in({
      m9_inst_col_repair_in[12:6], c1_gate1_m9_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts39), .ren(ren_ts39), .async_rst(m9_inst_async_rst), .fastsleep(m9_inst_fastsleep), 
      .deepsleep(m9_inst_deepsleep), .sbc(m9_inst_sbc), .shutoff(m9_inst_shutoff), 
      .mce(m9_inst_mce), .stbyp(m9_inst_stbyp), .rmce(m9_inst_rmce), .wmce(m9_inst_wmce), 
      .wpulse(m9_inst_wpulse), .wa_disable(m9_inst_wa_disable), .wa(m9_inst_wa), 
      .ra(m9_inst_ra), .global_rrow_en_in(m9_inst_global_rrow_en_in), .isolation_control_in(m9_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m9_inst_dpslp_or_shutoffout), .shutoffout(m9_inst_shutoffout), 
      .adr(adr_ts39), .din(din_ts39), .q(m9_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m10_inst(
      .row_repair_in({m10_inst_row_repair_in[25:21], 
      c1_gate1_m10_bisr_inst_Q[15:8], m10_inst_row_repair_in[12:8], 
      c1_gate1_m10_bisr_inst_Q[7:0]}), .col_repair_in({
      m10_inst_col_repair_in[12:6], c1_gate1_m10_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen), .ren(ren), .async_rst(m10_inst_async_rst), .fastsleep(m10_inst_fastsleep), 
      .deepsleep(m10_inst_deepsleep), .sbc(m10_inst_sbc), .shutoff(m10_inst_shutoff), 
      .mce(m10_inst_mce), .stbyp(m10_inst_stbyp), .rmce(m10_inst_rmce), .wmce(m10_inst_wmce), 
      .wpulse(m10_inst_wpulse), .wa_disable(m10_inst_wa_disable), .wa(m10_inst_wa), 
      .ra(m10_inst_ra), .global_rrow_en_in(m10_inst_global_rrow_en_in), .isolation_control_in(m10_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m10_inst_dpslp_or_shutoffout), .shutoffout(m10_inst_shutoffout), 
      .adr(adr), .din(din), .q(m10_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m11_inst(
      .row_repair_in({m11_inst_row_repair_in[25:21], 
      c1_gate1_m11_bisr_inst_Q[15:8], m11_inst_row_repair_in[12:8], 
      c1_gate1_m11_bisr_inst_Q[7:0]}), .col_repair_in({
      m11_inst_col_repair_in[12:6], c1_gate1_m11_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts1), .ren(ren_ts1), .async_rst(m11_inst_async_rst), .fastsleep(m11_inst_fastsleep), 
      .deepsleep(m11_inst_deepsleep), .sbc(m11_inst_sbc), .shutoff(m11_inst_shutoff), 
      .mce(m11_inst_mce), .stbyp(m11_inst_stbyp), .rmce(m11_inst_rmce), .wmce(m11_inst_wmce), 
      .wpulse(m11_inst_wpulse), .wa_disable(m11_inst_wa_disable), .wa(m11_inst_wa), 
      .ra(m11_inst_ra), .global_rrow_en_in(m11_inst_global_rrow_en_in), .isolation_control_in(m11_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m11_inst_dpslp_or_shutoffout), .shutoffout(m11_inst_shutoffout), 
      .adr(adr_ts1), .din(din_ts1), .q(m11_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m12_inst(
      .row_repair_in({m12_inst_row_repair_in[25:21], 
      c1_gate1_m12_bisr_inst_Q[15:8], m12_inst_row_repair_in[12:8], 
      c1_gate1_m12_bisr_inst_Q[7:0]}), .col_repair_in({
      m12_inst_col_repair_in[12:6], c1_gate1_m12_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts2), .ren(ren_ts2), .async_rst(m12_inst_async_rst), .fastsleep(m12_inst_fastsleep), 
      .deepsleep(m12_inst_deepsleep), .sbc(m12_inst_sbc), .shutoff(m12_inst_shutoff), 
      .mce(m12_inst_mce), .stbyp(m12_inst_stbyp), .rmce(m12_inst_rmce), .wmce(m12_inst_wmce), 
      .wpulse(m12_inst_wpulse), .wa_disable(m12_inst_wa_disable), .wa(m12_inst_wa), 
      .ra(m12_inst_ra), .global_rrow_en_in(m12_inst_global_rrow_en_in), .isolation_control_in(m12_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m12_inst_dpslp_or_shutoffout), .shutoffout(m12_inst_shutoffout), 
      .adr(adr_ts2), .din(din_ts2), .q(m12_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m13_inst(
      .row_repair_in({m13_inst_row_repair_in[25:21], 
      c1_gate1_m13_bisr_inst_Q[15:8], m13_inst_row_repair_in[12:8], 
      c1_gate1_m13_bisr_inst_Q[7:0]}), .col_repair_in({
      m13_inst_col_repair_in[12:6], c1_gate1_m13_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts3), .ren(ren_ts3), .async_rst(m13_inst_async_rst), .fastsleep(m13_inst_fastsleep), 
      .deepsleep(m13_inst_deepsleep), .sbc(m13_inst_sbc), .shutoff(m13_inst_shutoff), 
      .mce(m13_inst_mce), .stbyp(m13_inst_stbyp), .rmce(m13_inst_rmce), .wmce(m13_inst_wmce), 
      .wpulse(m13_inst_wpulse), .wa_disable(m13_inst_wa_disable), .wa(m13_inst_wa), 
      .ra(m13_inst_ra), .global_rrow_en_in(m13_inst_global_rrow_en_in), .isolation_control_in(m13_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m13_inst_dpslp_or_shutoffout), .shutoffout(m13_inst_shutoffout), 
      .adr(adr_ts3), .din(din_ts3), .q(m13_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m14_inst(
      .row_repair_in({m14_inst_row_repair_in[25:21], 
      c1_gate1_m14_bisr_inst_Q[15:8], m14_inst_row_repair_in[12:8], 
      c1_gate1_m14_bisr_inst_Q[7:0]}), .col_repair_in({
      m14_inst_col_repair_in[12:6], c1_gate1_m14_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts4), .ren(ren_ts4), .async_rst(m14_inst_async_rst), .fastsleep(m14_inst_fastsleep), 
      .deepsleep(m14_inst_deepsleep), .sbc(m14_inst_sbc), .shutoff(m14_inst_shutoff), 
      .mce(m14_inst_mce), .stbyp(m14_inst_stbyp), .rmce(m14_inst_rmce), .wmce(m14_inst_wmce), 
      .wpulse(m14_inst_wpulse), .wa_disable(m14_inst_wa_disable), .wa(m14_inst_wa), 
      .ra(m14_inst_ra), .global_rrow_en_in(m14_inst_global_rrow_en_in), .isolation_control_in(m14_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m14_inst_dpslp_or_shutoffout), .shutoffout(m14_inst_shutoffout), 
      .adr(adr_ts4), .din(din_ts4), .q(m14_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m15_inst(
      .row_repair_in({m15_inst_row_repair_in[25:21], 
      c1_gate1_m15_bisr_inst_Q[15:8], m15_inst_row_repair_in[12:8], 
      c1_gate1_m15_bisr_inst_Q[7:0]}), .col_repair_in({
      m15_inst_col_repair_in[12:6], c1_gate1_m15_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts5), .ren(ren_ts5), .async_rst(m15_inst_async_rst), .fastsleep(m15_inst_fastsleep), 
      .deepsleep(m15_inst_deepsleep), .sbc(m15_inst_sbc), .shutoff(m15_inst_shutoff), 
      .mce(m15_inst_mce), .stbyp(m15_inst_stbyp), .rmce(m15_inst_rmce), .wmce(m15_inst_wmce), 
      .wpulse(m15_inst_wpulse), .wa_disable(m15_inst_wa_disable), .wa(m15_inst_wa), 
      .ra(m15_inst_ra), .global_rrow_en_in(m15_inst_global_rrow_en_in), .isolation_control_in(m15_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m15_inst_dpslp_or_shutoffout), .shutoffout(m15_inst_shutoffout), 
      .adr(adr_ts5), .din(din_ts5), .q(m15_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m16_inst(
      .row_repair_in({m16_inst_row_repair_in[25:21], 
      c1_gate1_m16_bisr_inst_Q[15:8], m16_inst_row_repair_in[12:8], 
      c1_gate1_m16_bisr_inst_Q[7:0]}), .col_repair_in({
      m16_inst_col_repair_in[12:6], c1_gate1_m16_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts6), .ren(ren_ts6), .async_rst(m16_inst_async_rst), .fastsleep(m16_inst_fastsleep), 
      .deepsleep(m16_inst_deepsleep), .sbc(m16_inst_sbc), .shutoff(m16_inst_shutoff), 
      .mce(m16_inst_mce), .stbyp(m16_inst_stbyp), .rmce(m16_inst_rmce), .wmce(m16_inst_wmce), 
      .wpulse(m16_inst_wpulse), .wa_disable(m16_inst_wa_disable), .wa(m16_inst_wa), 
      .ra(m16_inst_ra), .global_rrow_en_in(m16_inst_global_rrow_en_in), .isolation_control_in(m16_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m16_inst_dpslp_or_shutoffout), .shutoffout(m16_inst_shutoffout), 
      .adr(adr_ts6), .din(din_ts6), .q(m16_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m17_inst(
      .row_repair_in({m17_inst_row_repair_in[25:21], 
      c1_gate1_m17_bisr_inst_Q[15:8], m17_inst_row_repair_in[12:8], 
      c1_gate1_m17_bisr_inst_Q[7:0]}), .col_repair_in({
      m17_inst_col_repair_in[12:6], c1_gate1_m17_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts7), .ren(ren_ts7), .async_rst(m17_inst_async_rst), .fastsleep(m17_inst_fastsleep), 
      .deepsleep(m17_inst_deepsleep), .sbc(m17_inst_sbc), .shutoff(m17_inst_shutoff), 
      .mce(m17_inst_mce), .stbyp(m17_inst_stbyp), .rmce(m17_inst_rmce), .wmce(m17_inst_wmce), 
      .wpulse(m17_inst_wpulse), .wa_disable(m17_inst_wa_disable), .wa(m17_inst_wa), 
      .ra(m17_inst_ra), .global_rrow_en_in(m17_inst_global_rrow_en_in), .isolation_control_in(m17_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m17_inst_dpslp_or_shutoffout), .shutoffout(m17_inst_shutoffout), 
      .adr(adr_ts7), .din(din_ts7), .q(m17_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m18_inst(
      .row_repair_in({m18_inst_row_repair_in[25:21], 
      c1_gate1_m18_bisr_inst_Q[15:8], m18_inst_row_repair_in[12:8], 
      c1_gate1_m18_bisr_inst_Q[7:0]}), .col_repair_in({
      m18_inst_col_repair_in[12:6], c1_gate1_m18_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts8), .ren(ren_ts8), .async_rst(m18_inst_async_rst), .fastsleep(m18_inst_fastsleep), 
      .deepsleep(m18_inst_deepsleep), .sbc(m18_inst_sbc), .shutoff(m18_inst_shutoff), 
      .mce(m18_inst_mce), .stbyp(m18_inst_stbyp), .rmce(m18_inst_rmce), .wmce(m18_inst_wmce), 
      .wpulse(m18_inst_wpulse), .wa_disable(m18_inst_wa_disable), .wa(m18_inst_wa), 
      .ra(m18_inst_ra), .global_rrow_en_in(m18_inst_global_rrow_en_in), .isolation_control_in(m18_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m18_inst_dpslp_or_shutoffout), .shutoffout(m18_inst_shutoffout), 
      .adr(adr_ts8), .din(din_ts8), .q(m18_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m19_inst(
      .row_repair_in({m19_inst_row_repair_in[25:21], 
      c1_gate1_m19_bisr_inst_Q[15:8], m19_inst_row_repair_in[12:8], 
      c1_gate1_m19_bisr_inst_Q[7:0]}), .col_repair_in({
      m19_inst_col_repair_in[12:6], c1_gate1_m19_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts9), .ren(ren_ts9), .async_rst(m19_inst_async_rst), .fastsleep(m19_inst_fastsleep), 
      .deepsleep(m19_inst_deepsleep), .sbc(m19_inst_sbc), .shutoff(m19_inst_shutoff), 
      .mce(m19_inst_mce), .stbyp(m19_inst_stbyp), .rmce(m19_inst_rmce), .wmce(m19_inst_wmce), 
      .wpulse(m19_inst_wpulse), .wa_disable(m19_inst_wa_disable), .wa(m19_inst_wa), 
      .ra(m19_inst_ra), .global_rrow_en_in(m19_inst_global_rrow_en_in), .isolation_control_in(m19_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m19_inst_dpslp_or_shutoffout), .shutoffout(m19_inst_shutoffout), 
      .adr(adr_ts9), .din(din_ts9), .q(m19_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m20_inst(
      .row_repair_in({m20_inst_row_repair_in[25:21], 
      c1_gate1_m20_bisr_inst_Q[15:8], m20_inst_row_repair_in[12:8], 
      c1_gate1_m20_bisr_inst_Q[7:0]}), .col_repair_in({
      m20_inst_col_repair_in[12:6], c1_gate1_m20_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts11), .ren(ren_ts11), .async_rst(m20_inst_async_rst), .fastsleep(m20_inst_fastsleep), 
      .deepsleep(m20_inst_deepsleep), .sbc(m20_inst_sbc), .shutoff(m20_inst_shutoff), 
      .mce(m20_inst_mce), .stbyp(m20_inst_stbyp), .rmce(m20_inst_rmce), .wmce(m20_inst_wmce), 
      .wpulse(m20_inst_wpulse), .wa_disable(m20_inst_wa_disable), .wa(m20_inst_wa), 
      .ra(m20_inst_ra), .global_rrow_en_in(m20_inst_global_rrow_en_in), .isolation_control_in(m20_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m20_inst_dpslp_or_shutoffout), .shutoffout(m20_inst_shutoffout), 
      .adr(adr_ts11), .din(din_ts11), .q(m20_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m21_inst(
      .row_repair_in({m21_inst_row_repair_in[25:21], 
      c1_gate1_m21_bisr_inst_Q[15:8], m21_inst_row_repair_in[12:8], 
      c1_gate1_m21_bisr_inst_Q[7:0]}), .col_repair_in({
      m21_inst_col_repair_in[12:6], c1_gate1_m21_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts12), .ren(ren_ts12), .async_rst(m21_inst_async_rst), .fastsleep(m21_inst_fastsleep), 
      .deepsleep(m21_inst_deepsleep), .sbc(m21_inst_sbc), .shutoff(m21_inst_shutoff), 
      .mce(m21_inst_mce), .stbyp(m21_inst_stbyp), .rmce(m21_inst_rmce), .wmce(m21_inst_wmce), 
      .wpulse(m21_inst_wpulse), .wa_disable(m21_inst_wa_disable), .wa(m21_inst_wa), 
      .ra(m21_inst_ra), .global_rrow_en_in(m21_inst_global_rrow_en_in), .isolation_control_in(m21_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m21_inst_dpslp_or_shutoffout), .shutoffout(m21_inst_shutoffout), 
      .adr(adr_ts12), .din(din_ts12), .q(m21_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m22_inst(
      .row_repair_in({m22_inst_row_repair_in[25:21], 
      c1_gate1_m22_bisr_inst_Q[15:8], m22_inst_row_repair_in[12:8], 
      c1_gate1_m22_bisr_inst_Q[7:0]}), .col_repair_in({
      m22_inst_col_repair_in[12:6], c1_gate1_m22_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts13), .ren(ren_ts13), .async_rst(m22_inst_async_rst), .fastsleep(m22_inst_fastsleep), 
      .deepsleep(m22_inst_deepsleep), .sbc(m22_inst_sbc), .shutoff(m22_inst_shutoff), 
      .mce(m22_inst_mce), .stbyp(m22_inst_stbyp), .rmce(m22_inst_rmce), .wmce(m22_inst_wmce), 
      .wpulse(m22_inst_wpulse), .wa_disable(m22_inst_wa_disable), .wa(m22_inst_wa), 
      .ra(m22_inst_ra), .global_rrow_en_in(m22_inst_global_rrow_en_in), .isolation_control_in(m22_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m22_inst_dpslp_or_shutoffout), .shutoffout(m22_inst_shutoffout), 
      .adr(adr_ts13), .din(din_ts13), .q(m22_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m23_inst(
      .row_repair_in({m23_inst_row_repair_in[25:21], 
      c1_gate1_m23_bisr_inst_Q[15:8], m23_inst_row_repair_in[12:8], 
      c1_gate1_m23_bisr_inst_Q[7:0]}), .col_repair_in({
      m23_inst_col_repair_in[12:6], c1_gate1_m23_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts14), .ren(ren_ts14), .async_rst(m23_inst_async_rst), .fastsleep(m23_inst_fastsleep), 
      .deepsleep(m23_inst_deepsleep), .sbc(m23_inst_sbc), .shutoff(m23_inst_shutoff), 
      .mce(m23_inst_mce), .stbyp(m23_inst_stbyp), .rmce(m23_inst_rmce), .wmce(m23_inst_wmce), 
      .wpulse(m23_inst_wpulse), .wa_disable(m23_inst_wa_disable), .wa(m23_inst_wa), 
      .ra(m23_inst_ra), .global_rrow_en_in(m23_inst_global_rrow_en_in), .isolation_control_in(m23_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m23_inst_dpslp_or_shutoffout), .shutoffout(m23_inst_shutoffout), 
      .adr(adr_ts14), .din(din_ts14), .q(m23_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m24_inst(
      .row_repair_in({m24_inst_row_repair_in[25:21], 
      c1_gate1_m24_bisr_inst_Q[15:8], m24_inst_row_repair_in[12:8], 
      c1_gate1_m24_bisr_inst_Q[7:0]}), .col_repair_in({
      m24_inst_col_repair_in[12:6], c1_gate1_m24_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts15), .ren(ren_ts15), .async_rst(m24_inst_async_rst), .fastsleep(m24_inst_fastsleep), 
      .deepsleep(m24_inst_deepsleep), .sbc(m24_inst_sbc), .shutoff(m24_inst_shutoff), 
      .mce(m24_inst_mce), .stbyp(m24_inst_stbyp), .rmce(m24_inst_rmce), .wmce(m24_inst_wmce), 
      .wpulse(m24_inst_wpulse), .wa_disable(m24_inst_wa_disable), .wa(m24_inst_wa), 
      .ra(m24_inst_ra), .global_rrow_en_in(m24_inst_global_rrow_en_in), .isolation_control_in(m24_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m24_inst_dpslp_or_shutoffout), .shutoffout(m24_inst_shutoffout), 
      .adr(adr_ts15), .din(din_ts15), .q(m24_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m25_inst(
      .row_repair_in({m25_inst_row_repair_in[25:21], 
      c1_gate1_m25_bisr_inst_Q[15:8], m25_inst_row_repair_in[12:8], 
      c1_gate1_m25_bisr_inst_Q[7:0]}), .col_repair_in({
      m25_inst_col_repair_in[12:6], c1_gate1_m25_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts16), .ren(ren_ts16), .async_rst(m25_inst_async_rst), .fastsleep(m25_inst_fastsleep), 
      .deepsleep(m25_inst_deepsleep), .sbc(m25_inst_sbc), .shutoff(m25_inst_shutoff), 
      .mce(m25_inst_mce), .stbyp(m25_inst_stbyp), .rmce(m25_inst_rmce), .wmce(m25_inst_wmce), 
      .wpulse(m25_inst_wpulse), .wa_disable(m25_inst_wa_disable), .wa(m25_inst_wa), 
      .ra(m25_inst_ra), .global_rrow_en_in(m25_inst_global_rrow_en_in), .isolation_control_in(m25_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m25_inst_dpslp_or_shutoffout), .shutoffout(m25_inst_shutoffout), 
      .adr(adr_ts16), .din(din_ts16), .q(m25_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m26_inst(
      .row_repair_in({m26_inst_row_repair_in[25:21], 
      c1_gate1_m26_bisr_inst_Q[15:8], m26_inst_row_repair_in[12:8], 
      c1_gate1_m26_bisr_inst_Q[7:0]}), .col_repair_in({
      m26_inst_col_repair_in[12:6], c1_gate1_m26_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts17), .ren(ren_ts17), .async_rst(m26_inst_async_rst), .fastsleep(m26_inst_fastsleep), 
      .deepsleep(m26_inst_deepsleep), .sbc(m26_inst_sbc), .shutoff(m26_inst_shutoff), 
      .mce(m26_inst_mce), .stbyp(m26_inst_stbyp), .rmce(m26_inst_rmce), .wmce(m26_inst_wmce), 
      .wpulse(m26_inst_wpulse), .wa_disable(m26_inst_wa_disable), .wa(m26_inst_wa), 
      .ra(m26_inst_ra), .global_rrow_en_in(m26_inst_global_rrow_en_in), .isolation_control_in(m26_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m26_inst_dpslp_or_shutoffout), .shutoffout(m26_inst_shutoffout), 
      .adr(adr_ts17), .din(din_ts17), .q(m26_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m27_inst(
      .row_repair_in({m27_inst_row_repair_in[25:21], 
      c1_gate1_m27_bisr_inst_Q[15:8], m27_inst_row_repair_in[12:8], 
      c1_gate1_m27_bisr_inst_Q[7:0]}), .col_repair_in({
      m27_inst_col_repair_in[12:6], c1_gate1_m27_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts18), .ren(ren_ts18), .async_rst(m27_inst_async_rst), .fastsleep(m27_inst_fastsleep), 
      .deepsleep(m27_inst_deepsleep), .sbc(m27_inst_sbc), .shutoff(m27_inst_shutoff), 
      .mce(m27_inst_mce), .stbyp(m27_inst_stbyp), .rmce(m27_inst_rmce), .wmce(m27_inst_wmce), 
      .wpulse(m27_inst_wpulse), .wa_disable(m27_inst_wa_disable), .wa(m27_inst_wa), 
      .ra(m27_inst_ra), .global_rrow_en_in(m27_inst_global_rrow_en_in), .isolation_control_in(m27_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m27_inst_dpslp_or_shutoffout), .shutoffout(m27_inst_shutoffout), 
      .adr(adr_ts18), .din(din_ts18), .q(m27_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m28_inst(
      .row_repair_in({m28_inst_row_repair_in[25:21], 
      c1_gate1_m28_bisr_inst_Q[15:8], m28_inst_row_repair_in[12:8], 
      c1_gate1_m28_bisr_inst_Q[7:0]}), .col_repair_in({
      m28_inst_col_repair_in[12:6], c1_gate1_m28_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts19), .ren(ren_ts19), .async_rst(m28_inst_async_rst), .fastsleep(m28_inst_fastsleep), 
      .deepsleep(m28_inst_deepsleep), .sbc(m28_inst_sbc), .shutoff(m28_inst_shutoff), 
      .mce(m28_inst_mce), .stbyp(m28_inst_stbyp), .rmce(m28_inst_rmce), .wmce(m28_inst_wmce), 
      .wpulse(m28_inst_wpulse), .wa_disable(m28_inst_wa_disable), .wa(m28_inst_wa), 
      .ra(m28_inst_ra), .global_rrow_en_in(m28_inst_global_rrow_en_in), .isolation_control_in(m28_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m28_inst_dpslp_or_shutoffout), .shutoffout(m28_inst_shutoffout), 
      .adr(adr_ts19), .din(din_ts19), .q(m28_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m29_inst(
      .row_repair_in({m29_inst_row_repair_in[25:21], 
      c1_gate1_m29_bisr_inst_Q[15:8], m29_inst_row_repair_in[12:8], 
      c1_gate1_m29_bisr_inst_Q[7:0]}), .col_repair_in({
      m29_inst_col_repair_in[12:6], c1_gate1_m29_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts20), .ren(ren_ts20), .async_rst(m29_inst_async_rst), .fastsleep(m29_inst_fastsleep), 
      .deepsleep(m29_inst_deepsleep), .sbc(m29_inst_sbc), .shutoff(m29_inst_shutoff), 
      .mce(m29_inst_mce), .stbyp(m29_inst_stbyp), .rmce(m29_inst_rmce), .wmce(m29_inst_wmce), 
      .wpulse(m29_inst_wpulse), .wa_disable(m29_inst_wa_disable), .wa(m29_inst_wa), 
      .ra(m29_inst_ra), .global_rrow_en_in(m29_inst_global_rrow_en_in), .isolation_control_in(m29_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m29_inst_dpslp_or_shutoffout), .shutoffout(m29_inst_shutoffout), 
      .adr(adr_ts20), .din(din_ts20), .q(m29_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m30_inst(
      .row_repair_in({m30_inst_row_repair_in[25:21], 
      c1_gate1_m30_bisr_inst_Q[15:8], m30_inst_row_repair_in[12:8], 
      c1_gate1_m30_bisr_inst_Q[7:0]}), .col_repair_in({
      m30_inst_col_repair_in[12:6], c1_gate1_m30_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts22), .ren(ren_ts22), .async_rst(m30_inst_async_rst), .fastsleep(m30_inst_fastsleep), 
      .deepsleep(m30_inst_deepsleep), .sbc(m30_inst_sbc), .shutoff(m30_inst_shutoff), 
      .mce(m30_inst_mce), .stbyp(m30_inst_stbyp), .rmce(m30_inst_rmce), .wmce(m30_inst_wmce), 
      .wpulse(m30_inst_wpulse), .wa_disable(m30_inst_wa_disable), .wa(m30_inst_wa), 
      .ra(m30_inst_ra), .global_rrow_en_in(m30_inst_global_rrow_en_in), .isolation_control_in(m30_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m30_inst_dpslp_or_shutoffout), .shutoffout(m30_inst_shutoffout), 
      .adr(adr_ts22), .din(din_ts22), .q(m30_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m31_inst(
      .row_repair_in({m31_inst_row_repair_in[25:21], 
      c1_gate1_m31_bisr_inst_Q[15:8], m31_inst_row_repair_in[12:8], 
      c1_gate1_m31_bisr_inst_Q[7:0]}), .col_repair_in({
      m31_inst_col_repair_in[12:6], c1_gate1_m31_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts23), .ren(ren_ts23), .async_rst(m31_inst_async_rst), .fastsleep(m31_inst_fastsleep), 
      .deepsleep(m31_inst_deepsleep), .sbc(m31_inst_sbc), .shutoff(m31_inst_shutoff), 
      .mce(m31_inst_mce), .stbyp(m31_inst_stbyp), .rmce(m31_inst_rmce), .wmce(m31_inst_wmce), 
      .wpulse(m31_inst_wpulse), .wa_disable(m31_inst_wa_disable), .wa(m31_inst_wa), 
      .ra(m31_inst_ra), .global_rrow_en_in(m31_inst_global_rrow_en_in), .isolation_control_in(m31_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m31_inst_dpslp_or_shutoffout), .shutoffout(m31_inst_shutoffout), 
      .adr(adr_ts23), .din(din_ts23), .q(m31_inst_q_ts1)
  );
  ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper m32_inst(
      .row_repair_in({m32_inst_row_repair_in[25:21], 
      c1_gate1_m32_bisr_inst_Q[15:8], m32_inst_row_repair_in[12:8], 
      c1_gate1_m32_bisr_inst_Q[7:0]}), .col_repair_in({
      m32_inst_col_repair_in[12:6], c1_gate1_m32_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts24), .ren(ren_ts24), .async_rst(m32_inst_async_rst), .fastsleep(m32_inst_fastsleep), 
      .deepsleep(m32_inst_deepsleep), .sbc(m32_inst_sbc), .shutoff(m32_inst_shutoff), 
      .mce(m32_inst_mce), .stbyp(m32_inst_stbyp), .rmce(m32_inst_rmce), .wmce(m32_inst_wmce), 
      .wpulse(m32_inst_wpulse), .wa_disable(m32_inst_wa_disable), .wa(m32_inst_wa), 
      .ra(m32_inst_ra), .global_rrow_en_in(m32_inst_global_rrow_en_in), .isolation_control_in(m32_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m32_inst_dpslp_or_shutoffout), .shutoffout(m32_inst_shutoffout), 
      .adr(adr_ts24), .din(din_ts24), .q(m32_inst_q_ts1)
  );
  ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper m33_inst(
      .row_repair_in({m33_inst_row_repair_in[25:22], 
      c1_gate1_m33_bisr_inst_Q[17:9], m33_inst_row_repair_in[12:9], 
      c1_gate1_m33_bisr_inst_Q[8:0]}), .col_repair_in({
      m33_inst_col_repair_in[12:8], c1_gate1_m33_bisr_inst_Q[25:18]}), .clk(clk_clk_bbm), 
      .wen(wen_ts25), .ren(ren_ts25), .async_rst(m33_inst_async_rst), .fastsleep(m33_inst_fastsleep), 
      .deepsleep(m33_inst_deepsleep), .sbc(m33_inst_sbc), .shutoff(m33_inst_shutoff), 
      .mce(m33_inst_mce), .stbyp(m33_inst_stbyp), .rmce(m33_inst_rmce), .wmce(m33_inst_wmce), 
      .wpulse(m33_inst_wpulse), .wa_disable(m33_inst_wa_disable), .wa(m33_inst_wa), 
      .ra(m33_inst_ra), .global_rrow_en_in(m33_inst_global_rrow_en_in), .isolation_control_in(m33_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m33_inst_dpslp_or_shutoffout), .shutoffout(m33_inst_shutoffout), 
      .adr(adr_ts25), .din(din_ts25), .q(m33_inst_q_ts1)
  );
  ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper m34_inst(
      .row_repair_in({m34_inst_row_repair_in[25:22], 
      c1_gate1_m34_bisr_inst_Q[17:9], m34_inst_row_repair_in[12:9], 
      c1_gate1_m34_bisr_inst_Q[8:0]}), .col_repair_in({
      m34_inst_col_repair_in[12:8], c1_gate1_m34_bisr_inst_Q[25:18]}), .clk(clk_clk_bbm), 
      .wen(wen_ts26), .ren(ren_ts26), .async_rst(m34_inst_async_rst), .fastsleep(m34_inst_fastsleep), 
      .deepsleep(m34_inst_deepsleep), .sbc(m34_inst_sbc), .shutoff(m34_inst_shutoff), 
      .mce(m34_inst_mce), .stbyp(m34_inst_stbyp), .rmce(m34_inst_rmce), .wmce(m34_inst_wmce), 
      .wpulse(m34_inst_wpulse), .wa_disable(m34_inst_wa_disable), .wa(m34_inst_wa), 
      .ra(m34_inst_ra), .global_rrow_en_in(m34_inst_global_rrow_en_in), .isolation_control_in(m34_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m34_inst_dpslp_or_shutoffout), .shutoffout(m34_inst_shutoffout), 
      .adr(adr_ts26), .din(din_ts26), .q(m34_inst_q_ts1)
  );
  ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper m35_inst(
      .row_repair_in({m35_inst_row_repair_in[25:22], 
      c1_gate1_m35_bisr_inst_Q[17:9], m35_inst_row_repair_in[12:9], 
      c1_gate1_m35_bisr_inst_Q[8:0]}), .col_repair_in({
      m35_inst_col_repair_in[12:8], c1_gate1_m35_bisr_inst_Q[25:18]}), .clk(clk_clk_bbm), 
      .wen(wen_ts27), .ren(ren_ts27), .async_rst(m35_inst_async_rst), .fastsleep(m35_inst_fastsleep), 
      .deepsleep(m35_inst_deepsleep), .sbc(m35_inst_sbc), .shutoff(m35_inst_shutoff), 
      .mce(m35_inst_mce), .stbyp(m35_inst_stbyp), .rmce(m35_inst_rmce), .wmce(m35_inst_wmce), 
      .wpulse(m35_inst_wpulse), .wa_disable(m35_inst_wa_disable), .wa(m35_inst_wa), 
      .ra(m35_inst_ra), .global_rrow_en_in(m35_inst_global_rrow_en_in), .isolation_control_in(m35_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m35_inst_dpslp_or_shutoffout), .shutoffout(m35_inst_shutoffout), 
      .adr(adr_ts27), .din(din_ts27), .q(m35_inst_q_ts1)
  );
  ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper m36_inst(
      .row_repair_in({m36_inst_row_repair_in[25:22], 
      c1_gate1_m36_bisr_inst_Q[17:9], m36_inst_row_repair_in[12:9], 
      c1_gate1_m36_bisr_inst_Q[8:0]}), .col_repair_in({
      m36_inst_col_repair_in[12:8], c1_gate1_m36_bisr_inst_Q[25:18]}), .clk(clk_clk_bbm), 
      .wen(wen_ts28), .ren(ren_ts28), .async_rst(m36_inst_async_rst), .fastsleep(m36_inst_fastsleep), 
      .deepsleep(m36_inst_deepsleep), .sbc(m36_inst_sbc), .shutoff(m36_inst_shutoff), 
      .mce(m36_inst_mce), .stbyp(m36_inst_stbyp), .rmce(m36_inst_rmce), .wmce(m36_inst_wmce), 
      .wpulse(m36_inst_wpulse), .wa_disable(m36_inst_wa_disable), .wa(m36_inst_wa), 
      .ra(m36_inst_ra), .global_rrow_en_in(m36_inst_global_rrow_en_in), .isolation_control_in(m36_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m36_inst_dpslp_or_shutoffout), .shutoffout(m36_inst_shutoffout), 
      .adr(adr_ts28), .din(din_ts28), .q(m36_inst_q_ts1)
  );
  ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper m37_inst(
      .row_repair_in({m37_inst_row_repair_in[25:21], 
      c1_gate1_m37_bisr_inst_Q[15:8], m37_inst_row_repair_in[12:8], 
      c1_gate1_m37_bisr_inst_Q[7:0]}), .col_repair_in({
      m37_inst_col_repair_in[12:6], c1_gate1_m37_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts29), .ren(ren_ts29), .async_rst(m37_inst_async_rst), .fastsleep(m37_inst_fastsleep), 
      .deepsleep(m37_inst_deepsleep), .sbc(m37_inst_sbc), .shutoff(m37_inst_shutoff), 
      .mce(m37_inst_mce), .stbyp(m37_inst_stbyp), .rmce(m37_inst_rmce), .wmce(m37_inst_wmce), 
      .wpulse(m37_inst_wpulse), .wa_disable(m37_inst_wa_disable), .wa(m37_inst_wa), 
      .ra(m37_inst_ra), .global_rrow_en_in(m37_inst_global_rrow_en_in), .isolation_control_in(m37_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m37_inst_dpslp_or_shutoffout), .shutoffout(m37_inst_shutoffout), 
      .adr(adr_ts29), .din(din_ts29), .q(m37_inst_q_ts1)
  );
  ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper m38_inst(
      .row_repair_in({m38_inst_row_repair_in[25:21], 
      c1_gate1_m38_bisr_inst_Q[15:8], m38_inst_row_repair_in[12:8], 
      c1_gate1_m38_bisr_inst_Q[7:0]}), .col_repair_in({
      m38_inst_col_repair_in[12:6], c1_gate1_m38_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts30), .ren(ren_ts30), .async_rst(m38_inst_async_rst), .fastsleep(m38_inst_fastsleep), 
      .deepsleep(m38_inst_deepsleep), .sbc(m38_inst_sbc), .shutoff(m38_inst_shutoff), 
      .mce(m38_inst_mce), .stbyp(m38_inst_stbyp), .rmce(m38_inst_rmce), .wmce(m38_inst_wmce), 
      .wpulse(m38_inst_wpulse), .wa_disable(m38_inst_wa_disable), .wa(m38_inst_wa), 
      .ra(m38_inst_ra), .global_rrow_en_in(m38_inst_global_rrow_en_in), .isolation_control_in(m38_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m38_inst_dpslp_or_shutoffout), .shutoffout(m38_inst_shutoffout), 
      .adr(adr_ts30), .din(din_ts30), .q(m38_inst_q_ts1)
  );
  ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper m39_inst(
      .row_repair_in({m39_inst_row_repair_in[25:21], 
      c1_gate1_m39_bisr_inst_Q[15:8], m39_inst_row_repair_in[12:8], 
      c1_gate1_m39_bisr_inst_Q[7:0]}), .col_repair_in({
      m39_inst_col_repair_in[12:6], c1_gate1_m39_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts31), .ren(ren_ts31), .async_rst(m39_inst_async_rst), .fastsleep(m39_inst_fastsleep), 
      .deepsleep(m39_inst_deepsleep), .sbc(m39_inst_sbc), .shutoff(m39_inst_shutoff), 
      .mce(m39_inst_mce), .stbyp(m39_inst_stbyp), .rmce(m39_inst_rmce), .wmce(m39_inst_wmce), 
      .wpulse(m39_inst_wpulse), .wa_disable(m39_inst_wa_disable), .wa(m39_inst_wa), 
      .ra(m39_inst_ra), .global_rrow_en_in(m39_inst_global_rrow_en_in), .isolation_control_in(m39_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m39_inst_dpslp_or_shutoffout), .shutoffout(m39_inst_shutoffout), 
      .adr(adr_ts31), .din(din_ts31), .q(m39_inst_q_ts1)
  );
  ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper m40_inst(
      .row_repair_in({m40_inst_row_repair_in[25:21], 
      c1_gate1_m40_bisr_inst_Q[15:8], m40_inst_row_repair_in[12:8], 
      c1_gate1_m40_bisr_inst_Q[7:0]}), .col_repair_in({
      m40_inst_col_repair_in[12:6], c1_gate1_m40_bisr_inst_Q[21:16]}), .clk(clk_clk_bbm), 
      .wen(wen_ts33), .ren(ren_ts33), .async_rst(m40_inst_async_rst), .fastsleep(m40_inst_fastsleep), 
      .deepsleep(m40_inst_deepsleep), .sbc(m40_inst_sbc), .shutoff(m40_inst_shutoff), 
      .mce(m40_inst_mce), .stbyp(m40_inst_stbyp), .rmce(m40_inst_rmce), .wmce(m40_inst_wmce), 
      .wpulse(m40_inst_wpulse), .wa_disable(m40_inst_wa_disable), .wa(m40_inst_wa), 
      .ra(m40_inst_ra), .global_rrow_en_in(m40_inst_global_rrow_en_in), .isolation_control_in(m40_inst_isolation_control_in), 
      .dpslp_or_shutoffout(m40_inst_dpslp_or_shutoffout), .shutoffout(m40_inst_shutoffout), 
      .adr(adr_ts33), .din(din_ts33), .q(m40_inst_q_ts1)
  );
  firebird7_in_gate1_tessent_mbist_bap firebird7_in_gate1_tessent_mbist_bap_inst(
      .reset(reset), .ijtag_select(ijtag_select), .si(si), .capture_en(capture_en), 
      .shift_en(shift_en), .shift_en_R(), .update_en(update_en), .tck(tck), .to_interfaces_tck(to_interfaces_tck), 
      .to_controllers_tck(to_controllers_tck), .mcp_bounding_en(MCP_BOUNDING_EN), 
      .mcp_bounding_to_en(mcp_bounding_to_en), .scan_en(SCAN_SHIFT_EN), .scan_to_en(scan_to_en), 
      .memory_bypass_en(MEM_BYPASS_EN), .memory_bypass_to_en(memory_bypass_to_en), 
      .ltest_en(LV_TM), .ltest_to_en(ltest_to_en), .BIST_HOLD(BIST_HOLD), .ENABLE_MEM_RESET(ENABLE_MEM_RESET), 
      .REDUCED_ADDRESS_COUNT(REDUCED_ADDRESS_COUNT), .BIST_SELECT_TEST_DATA(BIST_SELECT_TEST_DATA), 
      .BIST_ALGO_MODE0(BIST_ALGO_MODE0), .BIST_ALGO_MODE1(BIST_ALGO_MODE1), .MEM_ARRAY_DUMP_MODE(MEM_ARRAY_DUMP_MODE), 
      .BIRA_EN(BIRA_EN), .BIST_DIAG_EN(BIST_DIAG_EN), .PRESERVE_FUSE_REGISTER(PRESERVE_FUSE_REGISTER), 
      .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), .BIST_ASYNC_RESET(BIST_ASYNC_RESET), 
      .FL_CNT_MODE0(FL_CNT_MODE0), .FL_CNT_MODE1(FL_CNT_MODE1), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .CHAIN_BYPASS_EN(), .TCK_MODE(), .BIST_SETUP({BIST_SETUP_ts2, 
      BIST_SETUP_ts1, BIST_SETUP}), .MBISTPG_GO(BIST_GO), .MBISTPG_DONE(BIST_DONE), 
      .bistEn(bistEn), .toBist(toBist), .fromBist(MBISTPG_SO), .so(so)
  );
  firebird7_in_gate1_tessent_mbist_c1_controller firebird7_in_gate1_tessent_mbist_c1_controller_inst(
      .MBIST_RA_PRSRV_FUSE_VAL(PRESERVE_FUSE_REGISTER), .MBISTPG_ALGO_SEL(7'b0000000), 
      .MBISTPG_ALGO_MODE({BIST_ALGO_MODE1, BIST_ALGO_MODE0}), .MBISTPG_MEM_RST(ENABLE_MEM_RESET), 
      .MBISTPG_REDUCED_ADDR_CNT_EN(REDUCED_ADDRESS_COUNT), .MEM_BYPASS_EN(memory_bypass_to_en), 
      .MCP_BOUNDING_EN(mcp_bounding_to_en), .MEM0_BIST_COLLAR_SO(BIST_SO_ts10), 
      .MEM1_BIST_COLLAR_SO(BIST_SO_ts21), .MEM2_BIST_COLLAR_SO(BIST_SO_ts32), .MEM3_BIST_COLLAR_SO(BIST_SO_ts34), 
      .MEM4_BIST_COLLAR_SO(BIST_SO_ts35), .MEM5_BIST_COLLAR_SO(BIST_SO_ts36), .MEM6_BIST_COLLAR_SO(BIST_SO_ts37), 
      .MEM7_BIST_COLLAR_SO(BIST_SO_ts38), .MEM8_BIST_COLLAR_SO(BIST_SO_ts39), .MEM9_BIST_COLLAR_SO(BIST_SO), 
      .MEM10_BIST_COLLAR_SO(BIST_SO_ts1), .MEM11_BIST_COLLAR_SO(BIST_SO_ts2), .MEM12_BIST_COLLAR_SO(BIST_SO_ts3), 
      .MEM13_BIST_COLLAR_SO(BIST_SO_ts4), .MEM14_BIST_COLLAR_SO(BIST_SO_ts5), .MEM15_BIST_COLLAR_SO(BIST_SO_ts6), 
      .MEM16_BIST_COLLAR_SO(BIST_SO_ts7), .MEM17_BIST_COLLAR_SO(BIST_SO_ts8), .MEM18_BIST_COLLAR_SO(BIST_SO_ts9), 
      .MEM19_BIST_COLLAR_SO(BIST_SO_ts11), .MEM20_BIST_COLLAR_SO(BIST_SO_ts12), 
      .MEM21_BIST_COLLAR_SO(BIST_SO_ts13), .MEM22_BIST_COLLAR_SO(BIST_SO_ts14), 
      .MEM23_BIST_COLLAR_SO(BIST_SO_ts15), .MEM24_BIST_COLLAR_SO(BIST_SO_ts16), 
      .MEM25_BIST_COLLAR_SO(BIST_SO_ts17), .MEM26_BIST_COLLAR_SO(BIST_SO_ts18), 
      .MEM27_BIST_COLLAR_SO(BIST_SO_ts19), .MEM28_BIST_COLLAR_SO(BIST_SO_ts20), 
      .MEM29_BIST_COLLAR_SO(BIST_SO_ts22), .MEM30_BIST_COLLAR_SO(BIST_SO_ts23), 
      .MEM31_BIST_COLLAR_SO(BIST_SO_ts24), .MEM32_BIST_COLLAR_SO(BIST_SO_ts25), 
      .MEM33_BIST_COLLAR_SO(BIST_SO_ts26), .MEM34_BIST_COLLAR_SO(BIST_SO_ts27), 
      .MEM35_BIST_COLLAR_SO(BIST_SO_ts28), .MEM36_BIST_COLLAR_SO(BIST_SO_ts29), 
      .MEM37_BIST_COLLAR_SO(BIST_SO_ts30), .MEM38_BIST_COLLAR_SO(BIST_SO_ts31), 
      .MEM39_BIST_COLLAR_SO(BIST_SO_ts33), .FL_CNT_MODE({FL_CNT_MODE1, 
      FL_CNT_MODE0}), .MBISTPG_BIRA_EN(BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_COLLAR_GO({BIST_GO_ts34, BIST_GO_ts32, BIST_GO_ts31, 
      BIST_GO_ts30, BIST_GO_ts29, BIST_GO_ts28, BIST_GO_ts27, BIST_GO_ts26, 
      BIST_GO_ts25, BIST_GO_ts24, BIST_GO_ts23, BIST_GO_ts21, BIST_GO_ts20, 
      BIST_GO_ts19, BIST_GO_ts18, BIST_GO_ts17, BIST_GO_ts16, BIST_GO_ts15, 
      BIST_GO_ts14, BIST_GO_ts13, BIST_GO_ts12, BIST_GO_ts10, BIST_GO_ts9, 
      BIST_GO_ts8, BIST_GO_ts7, BIST_GO_ts6, BIST_GO_ts5, BIST_GO_ts4, 
      BIST_GO_ts3, BIST_GO_ts2, BIST_GO_ts1, BIST_GO_ts40, BIST_GO_ts39, 
      BIST_GO_ts38, BIST_GO_ts37, BIST_GO_ts36, BIST_GO_ts35, BIST_GO_ts33, 
      BIST_GO_ts22, BIST_GO_ts11}), .MBISTPG_DIAG_EN(BIST_DIAG_EN), .BIST_CLK(clk_clk_bbm), 
      .BIST_SI(toBist), .BIST_HOLD(BIST_HOLD), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP({
      BIST_SETUP_ts1, BIST_SETUP}), .MBISTPG_TESTDATA_SELECT(BIST_SELECT_TEST_DATA), 
      .TCK(to_controllers_tck), .MBISTPG_EN(bistEn), .MBISTPG_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .LV_TM(ltest_to_en), .MBISTPG_MEM_ARRAY_DUMP_MODE(MEM_ARRAY_DUMP_MODE), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), 
      .MBISTPG_RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts7, BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, 
      BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .BIST_EXPECT_DATA({BIST_EXPECT_DATA_ts3, 
      BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, BIST_EXPECT_DATA}), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), 
      .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), .MEM0_BIST_COLLAR_SI(MEM0_BIST_COLLAR_SI), 
      .MEM1_BIST_COLLAR_SI(MEM1_BIST_COLLAR_SI), .MEM2_BIST_COLLAR_SI(MEM2_BIST_COLLAR_SI), 
      .MEM3_BIST_COLLAR_SI(MEM3_BIST_COLLAR_SI), .MEM4_BIST_COLLAR_SI(MEM4_BIST_COLLAR_SI), 
      .MEM5_BIST_COLLAR_SI(MEM5_BIST_COLLAR_SI), .MEM6_BIST_COLLAR_SI(MEM6_BIST_COLLAR_SI), 
      .MEM7_BIST_COLLAR_SI(MEM7_BIST_COLLAR_SI), .MEM8_BIST_COLLAR_SI(MEM8_BIST_COLLAR_SI), 
      .MEM9_BIST_COLLAR_SI(MEM9_BIST_COLLAR_SI), .MEM10_BIST_COLLAR_SI(MEM10_BIST_COLLAR_SI), 
      .MEM11_BIST_COLLAR_SI(MEM11_BIST_COLLAR_SI), .MEM12_BIST_COLLAR_SI(MEM12_BIST_COLLAR_SI), 
      .MEM13_BIST_COLLAR_SI(MEM13_BIST_COLLAR_SI), .MEM14_BIST_COLLAR_SI(MEM14_BIST_COLLAR_SI), 
      .MEM15_BIST_COLLAR_SI(MEM15_BIST_COLLAR_SI), .MEM16_BIST_COLLAR_SI(MEM16_BIST_COLLAR_SI), 
      .MEM17_BIST_COLLAR_SI(MEM17_BIST_COLLAR_SI), .MEM18_BIST_COLLAR_SI(MEM18_BIST_COLLAR_SI), 
      .MEM19_BIST_COLLAR_SI(MEM19_BIST_COLLAR_SI), .MEM20_BIST_COLLAR_SI(MEM20_BIST_COLLAR_SI), 
      .MEM21_BIST_COLLAR_SI(MEM21_BIST_COLLAR_SI), .MEM22_BIST_COLLAR_SI(MEM22_BIST_COLLAR_SI), 
      .MEM23_BIST_COLLAR_SI(MEM23_BIST_COLLAR_SI), .MEM24_BIST_COLLAR_SI(MEM24_BIST_COLLAR_SI), 
      .MEM25_BIST_COLLAR_SI(MEM25_BIST_COLLAR_SI), .MEM26_BIST_COLLAR_SI(MEM26_BIST_COLLAR_SI), 
      .MEM27_BIST_COLLAR_SI(MEM27_BIST_COLLAR_SI), .MEM28_BIST_COLLAR_SI(MEM28_BIST_COLLAR_SI), 
      .MEM29_BIST_COLLAR_SI(MEM29_BIST_COLLAR_SI), .MEM30_BIST_COLLAR_SI(MEM30_BIST_COLLAR_SI), 
      .MEM31_BIST_COLLAR_SI(MEM31_BIST_COLLAR_SI), .MEM32_BIST_COLLAR_SI(MEM32_BIST_COLLAR_SI), 
      .MEM33_BIST_COLLAR_SI(MEM33_BIST_COLLAR_SI), .MEM34_BIST_COLLAR_SI(MEM34_BIST_COLLAR_SI), 
      .MEM35_BIST_COLLAR_SI(MEM35_BIST_COLLAR_SI), .MEM36_BIST_COLLAR_SI(MEM36_BIST_COLLAR_SI), 
      .MEM37_BIST_COLLAR_SI(MEM37_BIST_COLLAR_SI), .MEM38_BIST_COLLAR_SI(MEM38_BIST_COLLAR_SI), 
      .MEM39_BIST_COLLAR_SI(MEM39_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), .BIST_COLLAR_DIAG_EN(BIST_COLLAR_DIAG_EN), 
      .BIST_COLLAR_BIRA_EN(BIST_COLLAR_BIRA_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .MBISTPG_SO(MBISTPG_SO), .PriorityColumn(PriorityColumn), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_CMP(BIST_CMP), 
      .BIST_COLLAR_EN0(BIST_COLLAR_EN0), .BIST_RUN_TO_COLLAR0(BIST_RUN_TO_COLLAR0), 
      .BIST_COLLAR_EN1(BIST_COLLAR_EN1), .BIST_RUN_TO_COLLAR1(BIST_RUN_TO_COLLAR1), 
      .BIST_COLLAR_EN2(BIST_COLLAR_EN2), .BIST_RUN_TO_COLLAR2(BIST_RUN_TO_COLLAR2), 
      .BIST_COLLAR_EN3(BIST_COLLAR_EN3), .BIST_RUN_TO_COLLAR3(BIST_RUN_TO_COLLAR3), 
      .BIST_COLLAR_EN4(BIST_COLLAR_EN4), .BIST_RUN_TO_COLLAR4(BIST_RUN_TO_COLLAR4), 
      .BIST_COLLAR_EN5(BIST_COLLAR_EN5), .BIST_RUN_TO_COLLAR5(BIST_RUN_TO_COLLAR5), 
      .BIST_COLLAR_EN6(BIST_COLLAR_EN6), .BIST_RUN_TO_COLLAR6(BIST_RUN_TO_COLLAR6), 
      .BIST_COLLAR_EN7(BIST_COLLAR_EN7), .BIST_RUN_TO_COLLAR7(BIST_RUN_TO_COLLAR7), 
      .BIST_COLLAR_EN8(BIST_COLLAR_EN8), .BIST_RUN_TO_COLLAR8(BIST_RUN_TO_COLLAR8), 
      .BIST_COLLAR_EN9(BIST_COLLAR_EN9), .BIST_RUN_TO_COLLAR9(BIST_RUN_TO_COLLAR9), 
      .BIST_COLLAR_EN10(BIST_COLLAR_EN10), .BIST_RUN_TO_COLLAR10(BIST_RUN_TO_COLLAR10), 
      .BIST_COLLAR_EN11(BIST_COLLAR_EN11), .BIST_RUN_TO_COLLAR11(BIST_RUN_TO_COLLAR11), 
      .BIST_COLLAR_EN12(BIST_COLLAR_EN12), .BIST_RUN_TO_COLLAR12(BIST_RUN_TO_COLLAR12), 
      .BIST_COLLAR_EN13(BIST_COLLAR_EN13), .BIST_RUN_TO_COLLAR13(BIST_RUN_TO_COLLAR13), 
      .BIST_COLLAR_EN14(BIST_COLLAR_EN14), .BIST_RUN_TO_COLLAR14(BIST_RUN_TO_COLLAR14), 
      .BIST_COLLAR_EN15(BIST_COLLAR_EN15), .BIST_RUN_TO_COLLAR15(BIST_RUN_TO_COLLAR15), 
      .BIST_COLLAR_EN16(BIST_COLLAR_EN16), .BIST_RUN_TO_COLLAR16(BIST_RUN_TO_COLLAR16), 
      .BIST_COLLAR_EN17(BIST_COLLAR_EN17), .BIST_RUN_TO_COLLAR17(BIST_RUN_TO_COLLAR17), 
      .BIST_COLLAR_EN18(BIST_COLLAR_EN18), .BIST_RUN_TO_COLLAR18(BIST_RUN_TO_COLLAR18), 
      .BIST_COLLAR_EN19(BIST_COLLAR_EN19), .BIST_RUN_TO_COLLAR19(BIST_RUN_TO_COLLAR19), 
      .BIST_COLLAR_EN20(BIST_COLLAR_EN20), .BIST_RUN_TO_COLLAR20(BIST_RUN_TO_COLLAR20), 
      .BIST_COLLAR_EN21(BIST_COLLAR_EN21), .BIST_RUN_TO_COLLAR21(BIST_RUN_TO_COLLAR21), 
      .BIST_COLLAR_EN22(BIST_COLLAR_EN22), .BIST_RUN_TO_COLLAR22(BIST_RUN_TO_COLLAR22), 
      .BIST_COLLAR_EN23(BIST_COLLAR_EN23), .BIST_RUN_TO_COLLAR23(BIST_RUN_TO_COLLAR23), 
      .BIST_COLLAR_EN24(BIST_COLLAR_EN24), .BIST_RUN_TO_COLLAR24(BIST_RUN_TO_COLLAR24), 
      .BIST_COLLAR_EN25(BIST_COLLAR_EN25), .BIST_RUN_TO_COLLAR25(BIST_RUN_TO_COLLAR25), 
      .BIST_COLLAR_EN26(BIST_COLLAR_EN26), .BIST_RUN_TO_COLLAR26(BIST_RUN_TO_COLLAR26), 
      .BIST_COLLAR_EN27(BIST_COLLAR_EN27), .BIST_RUN_TO_COLLAR27(BIST_RUN_TO_COLLAR27), 
      .BIST_COLLAR_EN28(BIST_COLLAR_EN28), .BIST_RUN_TO_COLLAR28(BIST_RUN_TO_COLLAR28), 
      .BIST_COLLAR_EN29(BIST_COLLAR_EN29), .BIST_RUN_TO_COLLAR29(BIST_RUN_TO_COLLAR29), 
      .BIST_COLLAR_EN30(BIST_COLLAR_EN30), .BIST_RUN_TO_COLLAR30(BIST_RUN_TO_COLLAR30), 
      .BIST_COLLAR_EN31(BIST_COLLAR_EN31), .BIST_RUN_TO_COLLAR31(BIST_RUN_TO_COLLAR31), 
      .BIST_COLLAR_EN32(BIST_COLLAR_EN32), .BIST_RUN_TO_COLLAR32(BIST_RUN_TO_COLLAR32), 
      .BIST_COLLAR_EN33(BIST_COLLAR_EN33), .BIST_RUN_TO_COLLAR33(BIST_RUN_TO_COLLAR33), 
      .BIST_COLLAR_EN34(BIST_COLLAR_EN34), .BIST_RUN_TO_COLLAR34(BIST_RUN_TO_COLLAR34), 
      .BIST_COLLAR_EN35(BIST_COLLAR_EN35), .BIST_RUN_TO_COLLAR35(BIST_RUN_TO_COLLAR35), 
      .BIST_COLLAR_EN36(BIST_COLLAR_EN36), .BIST_RUN_TO_COLLAR36(BIST_RUN_TO_COLLAR36), 
      .BIST_COLLAR_EN37(BIST_COLLAR_EN37), .BIST_RUN_TO_COLLAR37(BIST_RUN_TO_COLLAR37), 
      .BIST_COLLAR_EN38(BIST_COLLAR_EN38), .BIST_RUN_TO_COLLAR38(BIST_RUN_TO_COLLAR38), 
      .BIST_COLLAR_EN39(BIST_COLLAR_EN39), .BIST_RUN_TO_COLLAR39(BIST_RUN_TO_COLLAR39), 
      .CHKBCI_PHASE(CHKBCI_PHASE), .MBISTPG_GO(BIST_GO), .MBISTPG_STABLE(MBISTPG_STABLE), 
      .MBISTPG_DONE(BIST_DONE), .BIST_ON_TO_COLLAR(BIST_ON), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR)
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m1 m1_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m1_inst_wen), 
      .ren_IN(m1_inst_ren), .adr_IN(m1_inst_adr[9:0]), .din_IN(m1_inst_din[21:0]), 
      .q_IN(m1_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR0), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM0_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN0), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m1_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m1_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m1_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m1_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m1_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m1_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts10), .ren(ren_ts10), .adr(adr_ts10), .din(din_ts10), .q(m1_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts10), .BIST_GO(BIST_GO_ts11), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts10[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts10), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts10[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts10), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts10[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts10), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m2 m2_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m2_inst_wen), 
      .ren_IN(m2_inst_ren), .adr_IN(m2_inst_adr[9:0]), .din_IN(m2_inst_din[21:0]), 
      .q_IN(m2_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR1), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM1_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN1), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m2_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m2_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m2_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m2_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m2_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m2_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts21), .ren(ren_ts21), .adr(adr_ts21), .din(din_ts21), .q(m2_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts21), .BIST_GO(BIST_GO_ts22), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts21[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts21), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts21[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts21), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts21[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts21), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m3 m3_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m3_inst_wen), 
      .ren_IN(m3_inst_ren), .adr_IN(m3_inst_adr[9:0]), .din_IN(m3_inst_din[21:0]), 
      .q_IN(m3_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR2), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM2_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN2), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m3_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m3_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m3_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m3_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m3_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m3_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts32), .ren(ren_ts32), .adr(adr_ts32), .din(din_ts32), .q(m3_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts32), .BIST_GO(BIST_GO_ts33), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts32[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts32), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts32[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts32), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts32[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts32), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m4 m4_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m4_inst_wen), 
      .ren_IN(m4_inst_ren), .adr_IN(m4_inst_adr[9:0]), .din_IN(m4_inst_din[21:0]), 
      .q_IN(m4_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR3), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM3_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN3), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m4_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m4_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m4_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m4_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m4_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m4_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts34), .ren(ren_ts34), .adr(adr_ts34), .din(din_ts34), .q(m4_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts34), .BIST_GO(BIST_GO_ts35), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts34[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts34), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts34[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts34), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts34[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts34), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m5 m5_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m5_inst_wen), 
      .ren_IN(m5_inst_ren), .adr_IN(m5_inst_adr[9:0]), .din_IN(m5_inst_din[21:0]), 
      .q_IN(m5_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR4), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM4_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN4), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m5_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m5_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m5_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m5_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m5_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m5_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts35), .ren(ren_ts35), .adr(adr_ts35), .din(din_ts35), .q(m5_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts35), .BIST_GO(BIST_GO_ts36), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts35[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts35), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts35[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts35), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts35[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts35), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m6 m6_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m6_inst_wen), 
      .ren_IN(m6_inst_ren), .adr_IN(m6_inst_adr[9:0]), .din_IN(m6_inst_din[21:0]), 
      .q_IN(m6_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR5), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM5_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN5), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m6_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m6_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m6_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m6_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m6_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m6_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts36), .ren(ren_ts36), .adr(adr_ts36), .din(din_ts36), .q(m6_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts36), .BIST_GO(BIST_GO_ts37), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts36[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts36), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts36[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts36), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts36[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts36), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m7 m7_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m7_inst_wen), 
      .ren_IN(m7_inst_ren), .adr_IN(m7_inst_adr[9:0]), .din_IN(m7_inst_din[21:0]), 
      .q_IN(m7_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR6), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM6_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN6), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m7_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m7_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m7_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m7_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m7_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m7_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts37), .ren(ren_ts37), .adr(adr_ts37), .din(din_ts37), .q(m7_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts37), .BIST_GO(BIST_GO_ts38), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts37[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts37), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts37[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts37), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts37[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts37), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m8 m8_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m8_inst_wen), 
      .ren_IN(m8_inst_ren), .adr_IN(m8_inst_adr[9:0]), .din_IN(m8_inst_din[21:0]), 
      .q_IN(m8_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR7), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM7_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN7), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m8_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m8_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m8_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m8_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m8_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m8_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts38), .ren(ren_ts38), .adr(adr_ts38), .din(din_ts38), .q(m8_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts38), .BIST_GO(BIST_GO_ts39), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts38[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts38), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts38[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts38), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts38[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts38), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m9 m9_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m9_inst_wen), 
      .ren_IN(m9_inst_ren), .adr_IN(m9_inst_adr[9:0]), .din_IN(m9_inst_din[21:0]), 
      .q_IN(m9_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR8), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM8_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN8), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m9_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m9_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m9_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m9_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m9_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m9_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts39), .ren(ren_ts39), .adr(adr_ts39), .din(din_ts39), .q(m9_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts39), .BIST_GO(BIST_GO_ts40), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts39[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts39), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts39[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts39), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts39[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts39), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m10 m10_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m10_inst_wen), 
      .ren_IN(m10_inst_ren), .adr_IN(m10_inst_adr[9:0]), .din_IN(m10_inst_din[21:0]), 
      .q_IN(m10_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR9), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM9_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN9), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m10_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m10_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m10_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m10_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m10_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m10_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen), .ren(ren), .adr(adr), .din(din), .q(m10_inst_q[21:0]), .SCAN_OBS_FLOPS(), 
      .BIST_SO(BIST_SO), .BIST_GO(BIST_GO_ts1), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m11 m11_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m11_inst_wen), 
      .ren_IN(m11_inst_ren), .adr_IN(m11_inst_adr[9:0]), .din_IN(m11_inst_din[21:0]), 
      .q_IN(m11_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR10), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM10_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN10), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m11_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m11_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m11_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m11_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m11_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m11_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts1), .ren(ren_ts1), .adr(adr_ts1), .din(din_ts1), .q(m11_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts1), .BIST_GO(BIST_GO_ts2), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts1[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts1), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts1[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts1), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts1[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts1), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m12 m12_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m12_inst_wen), 
      .ren_IN(m12_inst_ren), .adr_IN(m12_inst_adr[9:0]), .din_IN(m12_inst_din[21:0]), 
      .q_IN(m12_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR11), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM11_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN11), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m12_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m12_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m12_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m12_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m12_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m12_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts2), .ren(ren_ts2), .adr(adr_ts2), .din(din_ts2), .q(m12_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts2), .BIST_GO(BIST_GO_ts3), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts2[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts2), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts2[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts2), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts2[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts2), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m13 m13_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m13_inst_wen), 
      .ren_IN(m13_inst_ren), .adr_IN(m13_inst_adr[9:0]), .din_IN(m13_inst_din[21:0]), 
      .q_IN(m13_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR12), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM12_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN12), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m13_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m13_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m13_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m13_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m13_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m13_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts3), .ren(ren_ts3), .adr(adr_ts3), .din(din_ts3), .q(m13_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts3), .BIST_GO(BIST_GO_ts4), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts3[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts3), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts3[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts3), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts3[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts3), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m14 m14_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m14_inst_wen), 
      .ren_IN(m14_inst_ren), .adr_IN(m14_inst_adr[9:0]), .din_IN(m14_inst_din[21:0]), 
      .q_IN(m14_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR13), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM13_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN13), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m14_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m14_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m14_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m14_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m14_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m14_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts4), .ren(ren_ts4), .adr(adr_ts4), .din(din_ts4), .q(m14_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts4), .BIST_GO(BIST_GO_ts5), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts4[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts4), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts4[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts4), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts4[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts4), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m15 m15_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m15_inst_wen), 
      .ren_IN(m15_inst_ren), .adr_IN(m15_inst_adr[9:0]), .din_IN(m15_inst_din[21:0]), 
      .q_IN(m15_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR14), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM14_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN14), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m15_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m15_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m15_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m15_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m15_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m15_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts5), .ren(ren_ts5), .adr(adr_ts5), .din(din_ts5), .q(m15_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts5), .BIST_GO(BIST_GO_ts6), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts5[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts5), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts5[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts5), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts5[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts5), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m16 m16_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m16_inst_wen), 
      .ren_IN(m16_inst_ren), .adr_IN(m16_inst_adr[9:0]), .din_IN(m16_inst_din[21:0]), 
      .q_IN(m16_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR15), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM15_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN15), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m16_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m16_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m16_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m16_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m16_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m16_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts6), .ren(ren_ts6), .adr(adr_ts6), .din(din_ts6), .q(m16_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts6), .BIST_GO(BIST_GO_ts7), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts6[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts6), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts6[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts6), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts6[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts6), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m17 m17_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m17_inst_wen), 
      .ren_IN(m17_inst_ren), .adr_IN(m17_inst_adr[9:0]), .din_IN(m17_inst_din[21:0]), 
      .q_IN(m17_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR16), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM16_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN16), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m17_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m17_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m17_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m17_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m17_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m17_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts7), .ren(ren_ts7), .adr(adr_ts7), .din(din_ts7), .q(m17_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts7), .BIST_GO(BIST_GO_ts8), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts7[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts7), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts7[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts7), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts7[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts7), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m18 m18_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m18_inst_wen), 
      .ren_IN(m18_inst_ren), .adr_IN(m18_inst_adr[9:0]), .din_IN(m18_inst_din[21:0]), 
      .q_IN(m18_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR17), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM17_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN17), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m18_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m18_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m18_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m18_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m18_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m18_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts8), .ren(ren_ts8), .adr(adr_ts8), .din(din_ts8), .q(m18_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts8), .BIST_GO(BIST_GO_ts9), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts8[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts8), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts8[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts8), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts8[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts8), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m19 m19_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m19_inst_wen), 
      .ren_IN(m19_inst_ren), .adr_IN(m19_inst_adr[9:0]), .din_IN(m19_inst_din[21:0]), 
      .q_IN(m19_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR18), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM18_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN18), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m19_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m19_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m19_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m19_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m19_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m19_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts9), .ren(ren_ts9), .adr(adr_ts9), .din(din_ts9), .q(m19_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts9), .BIST_GO(BIST_GO_ts10), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts9[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts9), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts9[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts9), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts9[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts9), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m20 m20_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m20_inst_wen), 
      .ren_IN(m20_inst_ren), .adr_IN(m20_inst_adr[9:0]), .din_IN(m20_inst_din[21:0]), 
      .q_IN(m20_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR19), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM19_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN19), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m20_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m20_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m20_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m20_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m20_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m20_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts11), .ren(ren_ts11), .adr(adr_ts11), .din(din_ts11), .q(m20_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts11), .BIST_GO(BIST_GO_ts12), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts11[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts11), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts11[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts11), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts11[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts11), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m21 m21_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m21_inst_wen), 
      .ren_IN(m21_inst_ren), .adr_IN(m21_inst_adr[9:0]), .din_IN(m21_inst_din[21:0]), 
      .q_IN(m21_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR20), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM20_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN20), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m21_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m21_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m21_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m21_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m21_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m21_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts12), .ren(ren_ts12), .adr(adr_ts12), .din(din_ts12), .q(m21_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts12), .BIST_GO(BIST_GO_ts13), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts12[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts12), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts12[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts12), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts12[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts12), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m22 m22_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m22_inst_wen), 
      .ren_IN(m22_inst_ren), .adr_IN(m22_inst_adr[9:0]), .din_IN(m22_inst_din[21:0]), 
      .q_IN(m22_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR21), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM21_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN21), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m22_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m22_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m22_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m22_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m22_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m22_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts13), .ren(ren_ts13), .adr(adr_ts13), .din(din_ts13), .q(m22_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts13), .BIST_GO(BIST_GO_ts14), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts13[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts13), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts13[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts13), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts13[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts13), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m23 m23_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m23_inst_wen), 
      .ren_IN(m23_inst_ren), .adr_IN(m23_inst_adr[9:0]), .din_IN(m23_inst_din[21:0]), 
      .q_IN(m23_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR22), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM22_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN22), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m23_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m23_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m23_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m23_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m23_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m23_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts14), .ren(ren_ts14), .adr(adr_ts14), .din(din_ts14), .q(m23_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts14), .BIST_GO(BIST_GO_ts15), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts14[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts14), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts14[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts14), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts14[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts14), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m24 m24_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m24_inst_wen), 
      .ren_IN(m24_inst_ren), .adr_IN(m24_inst_adr[9:0]), .din_IN(m24_inst_din[21:0]), 
      .q_IN(m24_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR23), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM23_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN23), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m24_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m24_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m24_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m24_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m24_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m24_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts15), .ren(ren_ts15), .adr(adr_ts15), .din(din_ts15), .q(m24_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts15), .BIST_GO(BIST_GO_ts16), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts15[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts15), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts15[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts15), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts15[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts15), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m25 m25_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m25_inst_wen), 
      .ren_IN(m25_inst_ren), .adr_IN(m25_inst_adr[9:0]), .din_IN(m25_inst_din[21:0]), 
      .q_IN(m25_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR24), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM24_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN24), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m25_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m25_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m25_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m25_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m25_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m25_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts16), .ren(ren_ts16), .adr(adr_ts16), .din(din_ts16), .q(m25_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts16), .BIST_GO(BIST_GO_ts17), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts16[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts16), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts16[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts16), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts16[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts16), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m26 m26_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m26_inst_wen), 
      .ren_IN(m26_inst_ren), .adr_IN(m26_inst_adr[9:0]), .din_IN(m26_inst_din[21:0]), 
      .q_IN(m26_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR25), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM25_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN25), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m26_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m26_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m26_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m26_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m26_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m26_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts17), .ren(ren_ts17), .adr(adr_ts17), .din(din_ts17), .q(m26_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts17), .BIST_GO(BIST_GO_ts18), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts17[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts17), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts17[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts17), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts17[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts17), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m27 m27_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m27_inst_wen), 
      .ren_IN(m27_inst_ren), .adr_IN(m27_inst_adr[9:0]), .din_IN(m27_inst_din[21:0]), 
      .q_IN(m27_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR26), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM26_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN26), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m27_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m27_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m27_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m27_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m27_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m27_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts18), .ren(ren_ts18), .adr(adr_ts18), .din(din_ts18), .q(m27_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts18), .BIST_GO(BIST_GO_ts19), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts18[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts18), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts18[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts18), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts18[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts18), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m28 m28_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m28_inst_wen), 
      .ren_IN(m28_inst_ren), .adr_IN(m28_inst_adr[9:0]), .din_IN(m28_inst_din[21:0]), 
      .q_IN(m28_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR27), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM27_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN27), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m28_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m28_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m28_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m28_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m28_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m28_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts19), .ren(ren_ts19), .adr(adr_ts19), .din(din_ts19), .q(m28_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts19), .BIST_GO(BIST_GO_ts20), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts19[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts19), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts19[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts19), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts19[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts19), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m29 m29_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m29_inst_wen), 
      .ren_IN(m29_inst_ren), .adr_IN(m29_inst_adr[9:0]), .din_IN(m29_inst_din[21:0]), 
      .q_IN(m29_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR28), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM28_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN28), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m29_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m29_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m29_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m29_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m29_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m29_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts20), .ren(ren_ts20), .adr(adr_ts20), .din(din_ts20), .q(m29_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts20), .BIST_GO(BIST_GO_ts21), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts20[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts20), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts20[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts20), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts20[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts20), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m30 m30_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m30_inst_wen), 
      .ren_IN(m30_inst_ren), .adr_IN(m30_inst_adr[9:0]), .din_IN(m30_inst_din[21:0]), 
      .q_IN(m30_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR29), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM29_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN29), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m30_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m30_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m30_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m30_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m30_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m30_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts22), .ren(ren_ts22), .adr(adr_ts22), .din(din_ts22), .q(m30_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts22), .BIST_GO(BIST_GO_ts23), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts22[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts22), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts22[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts22), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts22[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts22), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m31 m31_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m31_inst_wen), 
      .ren_IN(m31_inst_ren), .adr_IN(m31_inst_adr[9:0]), .din_IN(m31_inst_din[21:0]), 
      .q_IN(m31_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR30), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM30_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN30), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m31_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m31_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m31_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m31_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m31_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m31_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts23), .ren(ren_ts23), .adr(adr_ts23), .din(din_ts23), .q(m31_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts23), .BIST_GO(BIST_GO_ts24), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts23[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts23), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts23[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts23), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts23[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts23), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m32 m32_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m32_inst_wen), 
      .ren_IN(m32_inst_ren), .adr_IN(m32_inst_adr[9:0]), .din_IN(m32_inst_din[21:0]), 
      .q_IN(m32_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts2, BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR31), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM31_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN31), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m32_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m32_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m32_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m32_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m32_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m32_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts24), .ren(ren_ts24), .adr(adr_ts24), .din(din_ts24), .q(m32_inst_q[21:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts24), .BIST_GO(BIST_GO_ts25), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts24[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts24), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts24[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts24), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts24[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts24), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m33 m33_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m33_inst_wen), 
      .ren_IN(m33_inst_ren), .adr_IN(m33_inst_adr[9:0]), .din_IN(m33_inst_din[71:0]), 
      .q_IN(m33_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts7, 
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR32), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM32_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN32), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m33_bisr_inst_Q[8:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m33_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m33_bisr_inst_Q[17:10]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m33_bisr_inst_Q[9]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m33_bisr_inst_Q[25:19]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m33_bisr_inst_Q[18]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts25), .ren(ren_ts25), .adr(adr_ts25), .din(din_ts25), .q(m33_inst_q[71:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts25), .BIST_GO(BIST_GO_ts26), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts25[7:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts25), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts25[7:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts25), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts25[6:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts25), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m34 m34_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m34_inst_wen), 
      .ren_IN(m34_inst_ren), .adr_IN(m34_inst_adr[9:0]), .din_IN(m34_inst_din[71:0]), 
      .q_IN(m34_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts7, 
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR33), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM33_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN33), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m34_bisr_inst_Q[8:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m34_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m34_bisr_inst_Q[17:10]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m34_bisr_inst_Q[9]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m34_bisr_inst_Q[25:19]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m34_bisr_inst_Q[18]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts26), .ren(ren_ts26), .adr(adr_ts26), .din(din_ts26), .q(m34_inst_q[71:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts26), .BIST_GO(BIST_GO_ts27), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts26[7:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts26), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts26[7:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts26), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts26[6:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts26), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m35 m35_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m35_inst_wen), 
      .ren_IN(m35_inst_ren), .adr_IN(m35_inst_adr[9:0]), .din_IN(m35_inst_din[71:0]), 
      .q_IN(m35_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts7, 
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR34), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM34_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN34), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m35_bisr_inst_Q[8:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m35_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m35_bisr_inst_Q[17:10]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m35_bisr_inst_Q[9]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m35_bisr_inst_Q[25:19]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m35_bisr_inst_Q[18]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts27), .ren(ren_ts27), .adr(adr_ts27), .din(din_ts27), .q(m35_inst_q[71:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts27), .BIST_GO(BIST_GO_ts28), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts27[7:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts27), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts27[7:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts27), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts27[6:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts27), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m36 m36_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m36_inst_wen), 
      .ren_IN(m36_inst_ren), .adr_IN(m36_inst_adr[9:0]), .din_IN(m36_inst_din[71:0]), 
      .q_IN(m36_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts7, 
      BIST_ROW_ADD_ts6, BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, 
      BIST_ROW_ADD_ts2, BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({
      BIST_WRITE_DATA_ts3, BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, 
      BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), 
      .MEM_BYPASS_EN(memory_bypass_to_en), .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), 
      .BIST_ON(BIST_ON), .BIST_RUN(BIST_RUN_TO_COLLAR35), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), 
      .BIST_CLK(clk_clk_bbm), .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM35_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN35), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m36_bisr_inst_Q[8:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m36_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m36_bisr_inst_Q[17:10]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m36_bisr_inst_Q[9]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m36_bisr_inst_Q[25:19]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m36_bisr_inst_Q[18]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts28), .ren(ren_ts28), .adr(adr_ts28), .din(din_ts28), .q(m36_inst_q[71:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts28), .BIST_GO(BIST_GO_ts29), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts28[7:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts28), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts28[7:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts28), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts28[6:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts28), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m37 m37_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m37_inst_wen), 
      .ren_IN(m37_inst_ren), .adr_IN(m37_inst_adr[8:0]), .din_IN(m37_inst_din[31:0]), 
      .q_IN(m37_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts6, 
      BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts2, 
      BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({BIST_WRITE_DATA_ts3, 
      BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), 
      .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), .MEM_BYPASS_EN(memory_bypass_to_en), 
      .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), .BIST_ON(BIST_ON), 
      .BIST_RUN(BIST_RUN_TO_COLLAR36), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), .BIST_CLK(clk_clk_bbm), 
      .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM36_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN36), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m37_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m37_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m37_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m37_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m37_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m37_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts29), .ren(ren_ts29), .adr(adr_ts29), .din(din_ts29), .q(m37_inst_q[31:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts29), .BIST_GO(BIST_GO_ts30), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts29[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts29), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts29[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts29), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts29[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts29), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m38 m38_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m38_inst_wen), 
      .ren_IN(m38_inst_ren), .adr_IN(m38_inst_adr[8:0]), .din_IN(m38_inst_din[31:0]), 
      .q_IN(m38_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts6, 
      BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts2, 
      BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({BIST_WRITE_DATA_ts3, 
      BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), 
      .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), .MEM_BYPASS_EN(memory_bypass_to_en), 
      .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), .BIST_ON(BIST_ON), 
      .BIST_RUN(BIST_RUN_TO_COLLAR37), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), .BIST_CLK(clk_clk_bbm), 
      .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM37_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN37), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m38_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m38_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m38_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m38_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m38_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m38_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts30), .ren(ren_ts30), .adr(adr_ts30), .din(din_ts30), .q(m38_inst_q[31:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts30), .BIST_GO(BIST_GO_ts31), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts30[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts30), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts30[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts30), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts30[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts30), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m39 m39_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m39_inst_wen), 
      .ren_IN(m39_inst_ren), .adr_IN(m39_inst_adr[8:0]), .din_IN(m39_inst_din[31:0]), 
      .q_IN(m39_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts6, 
      BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts2, 
      BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({BIST_WRITE_DATA_ts3, 
      BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), 
      .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), .MEM_BYPASS_EN(memory_bypass_to_en), 
      .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), .BIST_ON(BIST_ON), 
      .BIST_RUN(BIST_RUN_TO_COLLAR38), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), .BIST_CLK(clk_clk_bbm), 
      .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM38_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN38), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m39_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m39_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m39_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m39_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m39_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m39_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts31), .ren(ren_ts31), .adr(adr_ts31), .din(din_ts31), .q(m39_inst_q[31:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts31), .BIST_GO(BIST_GO_ts32), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts31[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts31), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts31[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts31), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts31[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts31), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbist_c1_interface_m40 m40_interface_instance(
      .PriorityColumn(PriorityColumn), .BIST_CLEAR_BIRA(BIST_CLEAR_BIRA), .wen_IN(m40_inst_wen), 
      .ren_IN(m40_inst_ren), .adr_IN(m40_inst_adr[8:0]), .din_IN(m40_inst_din[31:0]), 
      .q_IN(m40_inst_q_ts1), .TCK(to_interfaces_tck), .BIST_CMP(BIST_CMP), .INCLUDE_MEM_RESULTS_REG(INCLUDE_MEM_RESULTS_REG), 
      .BIST_WRITEENABLE(BIST_WRITEENABLE), .BIST_READENABLE(BIST_READENABLE), .BIST_COL_ADD({
      BIST_COL_ADD_ts1, BIST_COL_ADD}), .BIST_ROW_ADD({BIST_ROW_ADD_ts6, 
      BIST_ROW_ADD_ts5, BIST_ROW_ADD_ts4, BIST_ROW_ADD_ts3, BIST_ROW_ADD_ts2, 
      BIST_ROW_ADD_ts1, BIST_ROW_ADD}), .BIST_WRITE_DATA({BIST_WRITE_DATA_ts3, 
      BIST_WRITE_DATA_ts2, BIST_WRITE_DATA_ts1, BIST_WRITE_DATA}), .CHKBCI_PHASE(CHKBCI_PHASE), 
      .BIST_TESTDATA_SELECT_TO_COLLAR(BIST_TESTDATA_SELECT_TO_COLLAR), .MEM_BYPASS_EN(memory_bypass_to_en), 
      .SCAN_SHIFT_EN(scan_to_en), .MCP_BOUNDING_EN(mcp_bounding_to_en), .BIST_ON(BIST_ON), 
      .BIST_RUN(BIST_RUN_TO_COLLAR39), .BIST_ASYNC_RESETN(BIST_ASYNC_RESET), .BIST_CLK(clk_clk_bbm), 
      .BIST_SHIFT_COLLAR(BIST_SHIFT_COLLAR), .BIST_EXPECT_DATA({
      BIST_EXPECT_DATA_ts3, BIST_EXPECT_DATA_ts2, BIST_EXPECT_DATA_ts1, 
      BIST_EXPECT_DATA}), .BIST_SI(MEM39_BIST_COLLAR_SI), .BIST_COLLAR_SETUP(BIST_COLLAR_SETUP), 
      .BIST_COLLAR_OPSET_SELECT(BIST_COLLAR_OPSET_SELECT), .BIST_COLLAR_HOLD(BIST_COLLAR_HOLD), 
      .BIST_BIRA_EN(BIST_COLLAR_BIRA_EN), .CHECK_REPAIR_NEEDED(CHECK_REPAIR_NEEDED), 
      .BIST_DIAG_EN(BIST_COLLAR_DIAG_EN), .BIST_CLEAR_DEFAULT(BIST_CLEAR_DEFAULT), 
      .BIST_CLEAR(BIST_CLEAR), .BIST_SETUP2(BIST_SETUP_ts2), .BIST_SETUP1(BIST_SETUP_ts1), 
      .BIST_SETUP0(BIST_SETUP), .LV_TM(ltest_to_en), .FREEZE_STOP_ERROR(FREEZE_STOP_ERROR), 
      .BIST_COLLAR_EN(BIST_COLLAR_EN39), .FROM_BISR_ALL_SROW0_FUSE_ADD_REG(c1_gate1_m40_bisr_inst_Q[7:1]), 
      .FROM_BISR_ALL_SROW0_ALLOC_REG(c1_gate1_m40_bisr_inst_Q[0]), .FROM_BISR_ALL_SROW1_FUSE_ADD_REG(c1_gate1_m40_bisr_inst_Q[15:9]), 
      .FROM_BISR_ALL_SROW1_ALLOC_REG(c1_gate1_m40_bisr_inst_Q[8]), .FROM_BISR_All_SCOL0_FUSE_REG(c1_gate1_m40_bisr_inst_Q[21:17]), 
      .FROM_BISR_All_SCOL0_ALLOC_REG(c1_gate1_m40_bisr_inst_Q[16]), .BIST_SHIFT_BIRA_COLLAR(BIST_SHIFT_BIRA_COLLAR), 
      .RESET_REG_SETUP2(MBISTPG_RESET_REG_SETUP2), .ERROR_CNT_ZERO(ERROR_CNT_ZERO), 
      .wen(wen_ts33), .ren(ren_ts33), .adr(adr_ts33), .din(din_ts33), .q(m40_inst_q[31:0]), 
      .SCAN_OBS_FLOPS(), .BIST_SO(BIST_SO_ts33), .BIST_GO(BIST_GO_ts34), .ALL_SROW0_FUSE_ADD_REG(ALL_SROW0_FUSE_ADD_REG_ts33[6:0]), 
      .ALL_SROW0_ALLOC_REG(ALL_SROW0_ALLOC_REG_ts33), .ALL_SROW1_FUSE_ADD_REG(ALL_SROW1_FUSE_ADD_REG_ts33[6:0]), 
      .ALL_SROW1_ALLOC_REG(ALL_SROW1_ALLOC_REG_ts33), .All_SCOL0_FUSE_REG(All_SCOL0_FUSE_REG_ts33[4:0]), 
      .All_SCOL0_ALLOC_REG(All_SCOL0_ALLOC_REG_ts33), .REPAIR_STATUS()
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m1_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(bisr_si), .SO(c1_gate1_m1_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts10[4:0], 
      All_SCOL0_ALLOC_REG_ts10, ALL_SROW1_FUSE_ADD_REG_ts10[6:0], 
      ALL_SROW1_ALLOC_REG_ts10, ALL_SROW0_FUSE_ADD_REG_ts10[6:0], 
      ALL_SROW0_ALLOC_REG_ts10}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m1_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m2_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m1_bisr_inst_SO), .SO(c1_gate1_m2_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts21[4:0], 
      All_SCOL0_ALLOC_REG_ts21, ALL_SROW1_FUSE_ADD_REG_ts21[6:0], 
      ALL_SROW1_ALLOC_REG_ts21, ALL_SROW0_FUSE_ADD_REG_ts21[6:0], 
      ALL_SROW0_ALLOC_REG_ts21}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m2_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m3_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m2_bisr_inst_SO), .SO(c1_gate1_m3_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts32[4:0], 
      All_SCOL0_ALLOC_REG_ts32, ALL_SROW1_FUSE_ADD_REG_ts32[6:0], 
      ALL_SROW1_ALLOC_REG_ts32, ALL_SROW0_FUSE_ADD_REG_ts32[6:0], 
      ALL_SROW0_ALLOC_REG_ts32}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m3_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m4_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m3_bisr_inst_SO), .SO(c1_gate1_m4_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts34[4:0], 
      All_SCOL0_ALLOC_REG_ts34, ALL_SROW1_FUSE_ADD_REG_ts34[6:0], 
      ALL_SROW1_ALLOC_REG_ts34, ALL_SROW0_FUSE_ADD_REG_ts34[6:0], 
      ALL_SROW0_ALLOC_REG_ts34}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m4_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m5_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m4_bisr_inst_SO), .SO(c1_gate1_m5_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts35[4:0], 
      All_SCOL0_ALLOC_REG_ts35, ALL_SROW1_FUSE_ADD_REG_ts35[6:0], 
      ALL_SROW1_ALLOC_REG_ts35, ALL_SROW0_FUSE_ADD_REG_ts35[6:0], 
      ALL_SROW0_ALLOC_REG_ts35}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m5_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m6_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m5_bisr_inst_SO), .SO(c1_gate1_m6_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts36[4:0], 
      All_SCOL0_ALLOC_REG_ts36, ALL_SROW1_FUSE_ADD_REG_ts36[6:0], 
      ALL_SROW1_ALLOC_REG_ts36, ALL_SROW0_FUSE_ADD_REG_ts36[6:0], 
      ALL_SROW0_ALLOC_REG_ts36}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m6_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m7_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m6_bisr_inst_SO), .SO(c1_gate1_m7_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts37[4:0], 
      All_SCOL0_ALLOC_REG_ts37, ALL_SROW1_FUSE_ADD_REG_ts37[6:0], 
      ALL_SROW1_ALLOC_REG_ts37, ALL_SROW0_FUSE_ADD_REG_ts37[6:0], 
      ALL_SROW0_ALLOC_REG_ts37}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m7_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m8_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m7_bisr_inst_SO), .SO(c1_gate1_m8_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts38[4:0], 
      All_SCOL0_ALLOC_REG_ts38, ALL_SROW1_FUSE_ADD_REG_ts38[6:0], 
      ALL_SROW1_ALLOC_REG_ts38, ALL_SROW0_FUSE_ADD_REG_ts38[6:0], 
      ALL_SROW0_ALLOC_REG_ts38}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m8_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m9_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m8_bisr_inst_SO), .SO(c1_gate1_m9_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts39[4:0], 
      All_SCOL0_ALLOC_REG_ts39, ALL_SROW1_FUSE_ADD_REG_ts39[6:0], 
      ALL_SROW1_ALLOC_REG_ts39, ALL_SROW0_FUSE_ADD_REG_ts39[6:0], 
      ALL_SROW0_ALLOC_REG_ts39}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m9_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m10_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m9_bisr_inst_SO), .SO(c1_gate1_m10_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG[4:0], All_SCOL0_ALLOC_REG, 
      ALL_SROW1_FUSE_ADD_REG[6:0], ALL_SROW1_ALLOC_REG, 
      ALL_SROW0_FUSE_ADD_REG[6:0], ALL_SROW0_ALLOC_REG}), .MSO(1'b0), .MSEL(1'b0), 
      .Q(c1_gate1_m10_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m11_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m10_bisr_inst_SO), .SO(c1_gate1_m11_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts1[4:0], 
      All_SCOL0_ALLOC_REG_ts1, ALL_SROW1_FUSE_ADD_REG_ts1[6:0], 
      ALL_SROW1_ALLOC_REG_ts1, ALL_SROW0_FUSE_ADD_REG_ts1[6:0], 
      ALL_SROW0_ALLOC_REG_ts1}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m11_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m12_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m11_bisr_inst_SO), .SO(c1_gate1_m12_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts2[4:0], 
      All_SCOL0_ALLOC_REG_ts2, ALL_SROW1_FUSE_ADD_REG_ts2[6:0], 
      ALL_SROW1_ALLOC_REG_ts2, ALL_SROW0_FUSE_ADD_REG_ts2[6:0], 
      ALL_SROW0_ALLOC_REG_ts2}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m12_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m13_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m12_bisr_inst_SO), .SO(c1_gate1_m13_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts3[4:0], 
      All_SCOL0_ALLOC_REG_ts3, ALL_SROW1_FUSE_ADD_REG_ts3[6:0], 
      ALL_SROW1_ALLOC_REG_ts3, ALL_SROW0_FUSE_ADD_REG_ts3[6:0], 
      ALL_SROW0_ALLOC_REG_ts3}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m13_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m14_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m13_bisr_inst_SO), .SO(c1_gate1_m14_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts4[4:0], 
      All_SCOL0_ALLOC_REG_ts4, ALL_SROW1_FUSE_ADD_REG_ts4[6:0], 
      ALL_SROW1_ALLOC_REG_ts4, ALL_SROW0_FUSE_ADD_REG_ts4[6:0], 
      ALL_SROW0_ALLOC_REG_ts4}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m14_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m15_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m14_bisr_inst_SO), .SO(c1_gate1_m15_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts5[4:0], 
      All_SCOL0_ALLOC_REG_ts5, ALL_SROW1_FUSE_ADD_REG_ts5[6:0], 
      ALL_SROW1_ALLOC_REG_ts5, ALL_SROW0_FUSE_ADD_REG_ts5[6:0], 
      ALL_SROW0_ALLOC_REG_ts5}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m15_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m16_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m15_bisr_inst_SO), .SO(c1_gate1_m16_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts6[4:0], 
      All_SCOL0_ALLOC_REG_ts6, ALL_SROW1_FUSE_ADD_REG_ts6[6:0], 
      ALL_SROW1_ALLOC_REG_ts6, ALL_SROW0_FUSE_ADD_REG_ts6[6:0], 
      ALL_SROW0_ALLOC_REG_ts6}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m16_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m17_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m16_bisr_inst_SO), .SO(c1_gate1_m17_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts7[4:0], 
      All_SCOL0_ALLOC_REG_ts7, ALL_SROW1_FUSE_ADD_REG_ts7[6:0], 
      ALL_SROW1_ALLOC_REG_ts7, ALL_SROW0_FUSE_ADD_REG_ts7[6:0], 
      ALL_SROW0_ALLOC_REG_ts7}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m17_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m18_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m17_bisr_inst_SO), .SO(c1_gate1_m18_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts8[4:0], 
      All_SCOL0_ALLOC_REG_ts8, ALL_SROW1_FUSE_ADD_REG_ts8[6:0], 
      ALL_SROW1_ALLOC_REG_ts8, ALL_SROW0_FUSE_ADD_REG_ts8[6:0], 
      ALL_SROW0_ALLOC_REG_ts8}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m18_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m19_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m18_bisr_inst_SO), .SO(c1_gate1_m19_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts9[4:0], 
      All_SCOL0_ALLOC_REG_ts9, ALL_SROW1_FUSE_ADD_REG_ts9[6:0], 
      ALL_SROW1_ALLOC_REG_ts9, ALL_SROW0_FUSE_ADD_REG_ts9[6:0], 
      ALL_SROW0_ALLOC_REG_ts9}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m19_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m20_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m19_bisr_inst_SO), .SO(c1_gate1_m20_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts11[4:0], 
      All_SCOL0_ALLOC_REG_ts11, ALL_SROW1_FUSE_ADD_REG_ts11[6:0], 
      ALL_SROW1_ALLOC_REG_ts11, ALL_SROW0_FUSE_ADD_REG_ts11[6:0], 
      ALL_SROW0_ALLOC_REG_ts11}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m20_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m21_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m20_bisr_inst_SO), .SO(c1_gate1_m21_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts12[4:0], 
      All_SCOL0_ALLOC_REG_ts12, ALL_SROW1_FUSE_ADD_REG_ts12[6:0], 
      ALL_SROW1_ALLOC_REG_ts12, ALL_SROW0_FUSE_ADD_REG_ts12[6:0], 
      ALL_SROW0_ALLOC_REG_ts12}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m21_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m22_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m21_bisr_inst_SO), .SO(c1_gate1_m22_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts13[4:0], 
      All_SCOL0_ALLOC_REG_ts13, ALL_SROW1_FUSE_ADD_REG_ts13[6:0], 
      ALL_SROW1_ALLOC_REG_ts13, ALL_SROW0_FUSE_ADD_REG_ts13[6:0], 
      ALL_SROW0_ALLOC_REG_ts13}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m22_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m23_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m22_bisr_inst_SO), .SO(c1_gate1_m23_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts14[4:0], 
      All_SCOL0_ALLOC_REG_ts14, ALL_SROW1_FUSE_ADD_REG_ts14[6:0], 
      ALL_SROW1_ALLOC_REG_ts14, ALL_SROW0_FUSE_ADD_REG_ts14[6:0], 
      ALL_SROW0_ALLOC_REG_ts14}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m23_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m24_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m23_bisr_inst_SO), .SO(c1_gate1_m24_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts15[4:0], 
      All_SCOL0_ALLOC_REG_ts15, ALL_SROW1_FUSE_ADD_REG_ts15[6:0], 
      ALL_SROW1_ALLOC_REG_ts15, ALL_SROW0_FUSE_ADD_REG_ts15[6:0], 
      ALL_SROW0_ALLOC_REG_ts15}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m24_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m25_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m24_bisr_inst_SO), .SO(c1_gate1_m25_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts16[4:0], 
      All_SCOL0_ALLOC_REG_ts16, ALL_SROW1_FUSE_ADD_REG_ts16[6:0], 
      ALL_SROW1_ALLOC_REG_ts16, ALL_SROW0_FUSE_ADD_REG_ts16[6:0], 
      ALL_SROW0_ALLOC_REG_ts16}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m25_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m26_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m25_bisr_inst_SO), .SO(c1_gate1_m26_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts17[4:0], 
      All_SCOL0_ALLOC_REG_ts17, ALL_SROW1_FUSE_ADD_REG_ts17[6:0], 
      ALL_SROW1_ALLOC_REG_ts17, ALL_SROW0_FUSE_ADD_REG_ts17[6:0], 
      ALL_SROW0_ALLOC_REG_ts17}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m26_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m27_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m26_bisr_inst_SO), .SO(c1_gate1_m27_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts18[4:0], 
      All_SCOL0_ALLOC_REG_ts18, ALL_SROW1_FUSE_ADD_REG_ts18[6:0], 
      ALL_SROW1_ALLOC_REG_ts18, ALL_SROW0_FUSE_ADD_REG_ts18[6:0], 
      ALL_SROW0_ALLOC_REG_ts18}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m27_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m28_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m27_bisr_inst_SO), .SO(c1_gate1_m28_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts19[4:0], 
      All_SCOL0_ALLOC_REG_ts19, ALL_SROW1_FUSE_ADD_REG_ts19[6:0], 
      ALL_SROW1_ALLOC_REG_ts19, ALL_SROW0_FUSE_ADD_REG_ts19[6:0], 
      ALL_SROW0_ALLOC_REG_ts19}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m28_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m29_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m28_bisr_inst_SO), .SO(c1_gate1_m29_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts20[4:0], 
      All_SCOL0_ALLOC_REG_ts20, ALL_SROW1_FUSE_ADD_REG_ts20[6:0], 
      ALL_SROW1_ALLOC_REG_ts20, ALL_SROW0_FUSE_ADD_REG_ts20[6:0], 
      ALL_SROW0_ALLOC_REG_ts20}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m29_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m30_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m29_bisr_inst_SO), .SO(c1_gate1_m30_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts22[4:0], 
      All_SCOL0_ALLOC_REG_ts22, ALL_SROW1_FUSE_ADD_REG_ts22[6:0], 
      ALL_SROW1_ALLOC_REG_ts22, ALL_SROW0_FUSE_ADD_REG_ts22[6:0], 
      ALL_SROW0_ALLOC_REG_ts22}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m30_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m31_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m30_bisr_inst_SO), .SO(c1_gate1_m31_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts23[4:0], 
      All_SCOL0_ALLOC_REG_ts23, ALL_SROW1_FUSE_ADD_REG_ts23[6:0], 
      ALL_SROW1_ALLOC_REG_ts23, ALL_SROW0_FUSE_ADD_REG_ts23[6:0], 
      ALL_SROW0_ALLOC_REG_ts23}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m31_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x22m8b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m32_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m31_bisr_inst_SO), .SO(c1_gate1_m32_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts24[4:0], 
      All_SCOL0_ALLOC_REG_ts24, ALL_SROW1_FUSE_ADD_REG_ts24[6:0], 
      ALL_SROW1_ALLOC_REG_ts24, ALL_SROW0_FUSE_ADD_REG_ts24[6:0], 
      ALL_SROW0_ALLOC_REG_ts24}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m32_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper c1_gate1_m33_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m32_bisr_inst_SO), .SO(c1_gate1_m33_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts25[6:0], 
      All_SCOL0_ALLOC_REG_ts25, ALL_SROW1_FUSE_ADD_REG_ts25[7:0], 
      ALL_SROW1_ALLOC_REG_ts25, ALL_SROW0_FUSE_ADD_REG_ts25[7:0], 
      ALL_SROW0_ALLOC_REG_ts25}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m33_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper c1_gate1_m34_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m33_bisr_inst_SO), .SO(c1_gate1_m34_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts26[6:0], 
      All_SCOL0_ALLOC_REG_ts26, ALL_SROW1_FUSE_ADD_REG_ts26[7:0], 
      ALL_SROW1_ALLOC_REG_ts26, ALL_SROW0_FUSE_ADD_REG_ts26[7:0], 
      ALL_SROW0_ALLOC_REG_ts26}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m34_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper c1_gate1_m35_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m34_bisr_inst_SO), .SO(c1_gate1_m35_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts27[6:0], 
      All_SCOL0_ALLOC_REG_ts27, ALL_SROW1_FUSE_ADD_REG_ts27[7:0], 
      ALL_SROW1_ALLOC_REG_ts27, ALL_SROW0_FUSE_ADD_REG_ts27[7:0], 
      ALL_SROW0_ALLOC_REG_ts27}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m35_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr1024x72m2b2s0c1r2p3d0a2_mem_wrapper c1_gate1_m36_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m35_bisr_inst_SO), .SO(c1_gate1_m36_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts28[6:0], 
      All_SCOL0_ALLOC_REG_ts28, ALL_SROW1_FUSE_ADD_REG_ts28[7:0], 
      ALL_SROW1_ALLOC_REG_ts28, ALL_SROW0_FUSE_ADD_REG_ts28[7:0], 
      ALL_SROW0_ALLOC_REG_ts28}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m36_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m37_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m36_bisr_inst_SO), .SO(c1_gate1_m37_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts29[4:0], 
      All_SCOL0_ALLOC_REG_ts29, ALL_SROW1_FUSE_ADD_REG_ts29[6:0], 
      ALL_SROW1_ALLOC_REG_ts29, ALL_SROW0_FUSE_ADD_REG_ts29[6:0], 
      ALL_SROW0_ALLOC_REG_ts29}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m37_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m38_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m37_bisr_inst_SO), .SO(c1_gate1_m38_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts30[4:0], 
      All_SCOL0_ALLOC_REG_ts30, ALL_SROW1_FUSE_ADD_REG_ts30[6:0], 
      ALL_SROW1_ALLOC_REG_ts30, ALL_SROW0_FUSE_ADD_REG_ts30[6:0], 
      ALL_SROW0_ALLOC_REG_ts30}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m38_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m39_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m38_bisr_inst_SO), .SO(c1_gate1_m39_bisr_inst_SO), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts31[4:0], 
      All_SCOL0_ALLOC_REG_ts31, ALL_SROW1_FUSE_ADD_REG_ts31[6:0], 
      ALL_SROW1_ALLOC_REG_ts31, ALL_SROW0_FUSE_ADD_REG_ts31[6:0], 
      ALL_SROW0_ALLOC_REG_ts31}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m39_bisr_inst_Q)
  );
  firebird7_in_gate1_tessent_mbisr_register_ip783hdspsr512x32m4b1s0c1r2p3d0a2_mem_wrapper c1_gate1_m40_bisr_inst(
      .CLK(bisr_clock), .RSTB(bisr_clear), .SI(c1_gate1_m39_bisr_inst_SO), .SO(bisr_so), 
      .SE(bisr_se), .D({All_SCOL0_FUSE_REG_ts33[4:0], 
      All_SCOL0_ALLOC_REG_ts33, ALL_SROW1_FUSE_ADD_REG_ts33[6:0], 
      ALL_SROW1_ALLOC_REG_ts33, ALL_SROW0_FUSE_ADD_REG_ts33[6:0], 
      ALL_SROW0_ALLOC_REG_ts33}), .MSO(1'b0), .MSEL(1'b0), .Q(c1_gate1_m40_bisr_inst_Q)
  );
endmodule

