//--------------------------------------------------------------------------------
//
//  Unpublished work. Copyright 2022 Siemens
//
//  This material contains trade secrets or otherwise confidential 
//  information owned by Siemens Industry Software Inc. or its affiliates 
//  (collectively, SISW), or its licensors. Access to and use of this 
//  information is strictly limited as set forth in the Customer's 
//  applicable agreements with SISW.
//
//--------------------------------------------------------------------------------
//  File created by: Tessent Shell
//          Version: 2022.4
//       Created on: Sun Oct 29 14:37:28 PDT 2023
//
//       IP version: 8
//--------------------------------------------------------------------------------


module firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_1 (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire [  3:0] edt_channels_in,
   output reg  [123:0] edt_scan_in,
   input  wire         from_next_segment,
   output wire         to_next_segment,
   output wire         unsegmented_bit_6
);
   reg    [ 14:0] lfsm_vec;
   reg    [ 14:0] lfsm_vec_lockup;

   // synopsys sync_set_reset edt_update
   always @(posedge edt_clock)
   begin : lfsm
      if (edt_update == 1'b1) begin
         lfsm_vec <= 15'b000000000000000;
      end
      else begin
         lfsm_vec[ 0] <= lfsm_vec[ 1] ^ edt_channels_in[1];
         lfsm_vec[ 1] <= lfsm_vec[ 2];
         lfsm_vec[ 2] <= lfsm_vec[ 3] ^ edt_channels_in[2];
         lfsm_vec[ 3] <= lfsm_vec[ 4];
         lfsm_vec[ 4] <= lfsm_vec[ 5] ^ edt_channels_in[3];
         lfsm_vec[ 5] <= lfsm_vec[ 6];
         lfsm_vec[ 6] <= lfsm_vec[ 7] ^ edt_channels_in[0];
         lfsm_vec[ 7] <= from_next_segment;
         lfsm_vec[ 8] <= lfsm_vec[ 9];
         lfsm_vec[ 9] <= lfsm_vec[10] ^ edt_channels_in[0];
         lfsm_vec[10] <= lfsm_vec[11] ^ lfsm_vec[ 4];
         lfsm_vec[11] <= lfsm_vec[12] ^ edt_channels_in[2];
         lfsm_vec[12] <= lfsm_vec[13];
         lfsm_vec[13] <= lfsm_vec[14] ^ edt_channels_in[3];
         lfsm_vec[14] <= lfsm_vec[ 0];
      end
   end

   assign to_next_segment    = lfsm_vec[ 8];
   assign unsegmented_bit_6  = lfsm_vec[ 6];

   always @(negedge edt_clock)
   begin : lockup_cells
      lfsm_vec_lockup <= lfsm_vec;
   end

   always @(lfsm_vec_lockup)
   begin : phase_shifter
      edt_scan_in[  0] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[  1] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[13];
      edt_scan_in[  2] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[  3] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[  4] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11];
      edt_scan_in[  5] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[  6] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[14];
      edt_scan_in[  7] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[  8] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[14];
      edt_scan_in[  9] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 10] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 11] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 12] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 13] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 14] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 15] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6];
      edt_scan_in[ 16] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 17] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 18] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 19] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 20] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 21] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 22] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 23] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 24] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 25] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 26] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 27] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 28] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 29] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 30] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 31] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 32] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[13] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 33] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 34] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 35] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 36] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 37] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 38] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 39] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 40] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 41] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 42] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 43] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 44] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 45] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 46] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 47] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 48] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4];
      edt_scan_in[ 49] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 50] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 51] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 52] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 53] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 54] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 55] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 5];
      edt_scan_in[ 56] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 57] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 58] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 59] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 60] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 61] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 62] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 63] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 64] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 65] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 66] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 67] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 68] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 69] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 70] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 71] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 72] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 73] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 74] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 75] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 76] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 77] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 78] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 79] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 80] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 81] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 82] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 83] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 84] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 85] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 86] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 87] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 88] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 89] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 90] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 91] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 92] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 93] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 94] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 95] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 96] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[14];
      edt_scan_in[ 97] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 98] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 99] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[14];
      edt_scan_in[100] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[101] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[102] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[103] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[104] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[14];
      edt_scan_in[105] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[106] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[107] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[108] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[14];
      edt_scan_in[109] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[110] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[111] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[112] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[113] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[114] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[115] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[116] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[117] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[118] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[14];
      edt_scan_in[119] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[120] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[14];
      edt_scan_in[121] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[122] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[123] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
   end

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_2 (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire [  3:0] edt_channels_in,
   output reg  [123:0] edt_scan_in,
   input  wire         from_previous_segment,
   output wire         to_previous_segment,
   input  wire         from_next_segment,
   output wire         to_next_segment,
   input  wire         unsegmented_bit_6
);
   reg    [ 13:0] lfsm_vec;
   reg    [ 13:0] lfsm_vec_lockup;

   // synopsys sync_set_reset edt_update
   always @(posedge edt_clock)
   begin : lfsm
      if (edt_update == 1'b1) begin
         lfsm_vec <= 14'b00000000000000;
      end
      else begin
         lfsm_vec[ 0] <= lfsm_vec[ 1];
         lfsm_vec[ 1] <= lfsm_vec[ 2];
         lfsm_vec[ 2] <= lfsm_vec[ 3] ^ edt_channels_in[2];
         lfsm_vec[ 3] <= lfsm_vec[ 4];
         lfsm_vec[ 4] <= lfsm_vec[ 5] ^ edt_channels_in[0];
         lfsm_vec[ 5] <= from_next_segment;
         lfsm_vec[ 6] <= lfsm_vec[ 7];
         lfsm_vec[ 7] <= lfsm_vec[ 8];
         lfsm_vec[ 8] <= lfsm_vec[ 9] ^ lfsm_vec[ 2];
         lfsm_vec[ 9] <= lfsm_vec[10] ^ edt_channels_in[3];
         lfsm_vec[10] <= lfsm_vec[11];
         lfsm_vec[11] <= lfsm_vec[12] ^ edt_channels_in[1];
         lfsm_vec[12] <= lfsm_vec[13] ^ unsegmented_bit_6;
         lfsm_vec[13] <= from_previous_segment ^ edt_channels_in[1];
      end
   end

   assign to_previous_segment = lfsm_vec[ 0];
   assign to_next_segment     = lfsm_vec[ 6];

   always @(negedge edt_clock)
   begin : lockup_cells
      lfsm_vec_lockup <= lfsm_vec;
   end

   always @(lfsm_vec_lockup)
   begin : phase_shifter
      edt_scan_in[  0] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[  1] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[  2] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[  3] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[  4] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[  5] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[  6] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[  7] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10];
      edt_scan_in[  8] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[  9] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 10] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 11] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 12] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 13] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 14] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 15] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6];
      edt_scan_in[ 16] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 17] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 18] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 19] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 20] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 21] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 22] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 23] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 24] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 25] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 26] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 27] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 28] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 29] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 30] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6];
      edt_scan_in[ 31] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 32] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 33] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 34] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 35] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 36] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 37] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 38] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 39] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 40] = lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 41] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 42] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 43] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 44] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 45] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 46] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 47] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 48] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 49] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 50] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 51] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 52] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 53] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 54] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 55] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 56] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 57] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 58] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 59] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 60] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 61] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 62] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 63] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 64] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 65] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 66] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 67] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 68] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 69] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 70] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 71] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 72] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 73] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 74] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 75] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 76] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 77] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 78] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 79] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 80] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10];
      edt_scan_in[ 81] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7];
      edt_scan_in[ 82] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 83] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 84] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 85] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 86] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6];
      edt_scan_in[ 87] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 88] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 89] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 90] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 91] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 92] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 93] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 94] = lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 95] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[ 96] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 97] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[ 98] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 99] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6];
      edt_scan_in[100] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[101] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[13];
      edt_scan_in[102] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[103] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11];
      edt_scan_in[104] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[105] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[106] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[107] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[108] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[109] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10];
      edt_scan_in[110] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[111] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[112] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11];
      edt_scan_in[113] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[114] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10];
      edt_scan_in[115] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[13];
      edt_scan_in[116] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[117] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[118] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10];
      edt_scan_in[119] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8];
      edt_scan_in[120] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[121] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10];
      edt_scan_in[122] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9];
      edt_scan_in[123] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6];
   end

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_3 (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire [  3:0] edt_channels_in,
   output reg  [122:0] edt_scan_in,
   input  wire         from_previous_segment,
   output wire         to_previous_segment
);
   reg    [ 13:0] lfsm_vec;
   reg    [ 13:0] lfsm_vec_lockup;

   // synopsys sync_set_reset edt_update
   always @(posedge edt_clock)
   begin : lfsm
      if (edt_update == 1'b1) begin
         lfsm_vec <= 14'b00000000000000;
      end
      else begin
         lfsm_vec[ 0] <= lfsm_vec[ 1];
         lfsm_vec[ 1] <= lfsm_vec[ 2];
         lfsm_vec[ 2] <= lfsm_vec[ 3];
         lfsm_vec[ 3] <= lfsm_vec[ 4];
         lfsm_vec[ 4] <= lfsm_vec[ 5];
         lfsm_vec[ 5] <= lfsm_vec[ 6] ^ edt_channels_in[3];
         lfsm_vec[ 6] <= lfsm_vec[ 7];
         lfsm_vec[ 7] <= lfsm_vec[ 8] ^ edt_channels_in[0];
         lfsm_vec[ 8] <= lfsm_vec[ 9];
         lfsm_vec[ 9] <= lfsm_vec[10] ^ edt_channels_in[1];
         lfsm_vec[10] <= lfsm_vec[11] ^ lfsm_vec[ 5];
         lfsm_vec[11] <= lfsm_vec[12] ^ edt_channels_in[2];
         lfsm_vec[12] <= lfsm_vec[13];
         lfsm_vec[13] <= from_previous_segment ^ lfsm_vec[ 1];
      end
   end

   assign to_previous_segment = lfsm_vec[ 0];

   always @(negedge edt_clock)
   begin : lockup_cells
      lfsm_vec_lockup <= lfsm_vec;
   end

   always @(lfsm_vec_lockup)
   begin : phase_shifter
      edt_scan_in[  0] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[  1] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[  2] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[  3] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[  4] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11];
      edt_scan_in[  5] = lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[  6] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[  7] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[  8] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[  9] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 10] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 11] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 12] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 13] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 14] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 15] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 16] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 17] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 18] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 19] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 20] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 21] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 22] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 23] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 24] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 25] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 26] = lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 27] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 28] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 29] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 30] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 31] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 32] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 33] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 34] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 35] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 36] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 37] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 38] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 39] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 40] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 41] = lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 42] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 43] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 44] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 45] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 46] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 47] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 48] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 49] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 50] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 51] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 52] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 53] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 54] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 55] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 56] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 57] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 58] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 59] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 60] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 61] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 62] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 63] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 64] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 65] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 66] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 67] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 68] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 69] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 70] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 71] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 72] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 73] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 74] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 75] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 76] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 77] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 78] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 79] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 80] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 81] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 82] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 83] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 84] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 85] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 86] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 87] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 88] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 89] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 90] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 91] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 92] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 93] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 94] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 95] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 96] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[11];
      edt_scan_in[ 97] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[ 98] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[ 99] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[12];
      edt_scan_in[100] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[13];
      edt_scan_in[101] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[102] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[103] = lfsm_vec_lockup[ 1] ^ lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[12];
      edt_scan_in[104] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[105] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[11];
      edt_scan_in[106] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[107] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[108] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
      edt_scan_in[109] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[110] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12];
      edt_scan_in[111] = lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[13];
      edt_scan_in[112] = lfsm_vec_lockup[ 6] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[113] = lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[114] = lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[11] ^ lfsm_vec_lockup[12];
      edt_scan_in[115] = lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[13];
      edt_scan_in[116] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 9] ^ lfsm_vec_lockup[13];
      edt_scan_in[117] = lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[12];
      edt_scan_in[118] = lfsm_vec_lockup[ 4] ^ lfsm_vec_lockup[ 7] ^ lfsm_vec_lockup[13];
      edt_scan_in[119] = lfsm_vec_lockup[ 0] ^ lfsm_vec_lockup[ 5] ^ lfsm_vec_lockup[11];
      edt_scan_in[120] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[12] ^ lfsm_vec_lockup[13];
      edt_scan_in[121] = lfsm_vec_lockup[ 2] ^ lfsm_vec_lockup[ 3] ^ lfsm_vec_lockup[13];
      edt_scan_in[122] = lfsm_vec_lockup[ 8] ^ lfsm_vec_lockup[10] ^ lfsm_vec_lockup[13];
   end

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_decompressor (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire [  3:0] edt_channels_in,
   output wire [370:0] edt_scan_in
);
   wire           seg_1to2;
   wire           seg_2to1;
   wire           seg_2to3;
   wire           seg_3to2;
   wire           unsegmented_bit_6;

   firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_1 segment1 (
      .edt_clock(edt_clock),
      .edt_update(edt_update),
      .edt_channels_in(edt_channels_in[3:0]),
      .edt_scan_in(edt_scan_in[123:0]),
      .from_next_segment(seg_2to1),
      .to_next_segment(seg_1to2),
      .unsegmented_bit_6(unsegmented_bit_6));
   firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_2 segment2 (
      .edt_clock(edt_clock),
      .edt_update(edt_update),
      .edt_channels_in(edt_channels_in[3:0]),
      .edt_scan_in(edt_scan_in[247:124]),
      .from_previous_segment(seg_1to2),
      .to_previous_segment(seg_2to1),
      .from_next_segment(seg_3to2),
      .to_next_segment(seg_2to3),
      .unsegmented_bit_6(unsegmented_bit_6));
   firebird7_in_gate2_tessent_edt_intest_edt_decompressor_segment_3 segment3 (
      .edt_clock(edt_clock),
      .edt_update(edt_update),
      .edt_channels_in(edt_channels_in[3:0]),
      .edt_scan_in(edt_scan_in[370:248]),
      .from_previous_segment(seg_2to3),
      .to_previous_segment(seg_3to2));
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_low_power_shift_decoder (
   input  wire [370:0] encoded_control,
   output wire [370:0] decoded_control
);
   assign decoded_control[  0] = encoded_control[  0];
   assign decoded_control[  1] = encoded_control[  1];
   assign decoded_control[  2] = encoded_control[  2];
   assign decoded_control[  3] = encoded_control[  3];
   assign decoded_control[  4] = encoded_control[  4];
   assign decoded_control[  5] = encoded_control[  5];
   assign decoded_control[  6] = encoded_control[  6];
   assign decoded_control[  7] = encoded_control[  7];
   assign decoded_control[  8] = encoded_control[  8];
   assign decoded_control[  9] = encoded_control[  9];
   assign decoded_control[ 10] = encoded_control[ 10];
   assign decoded_control[ 11] = encoded_control[ 11];
   assign decoded_control[ 12] = encoded_control[ 12];
   assign decoded_control[ 13] = encoded_control[ 13];
   assign decoded_control[ 14] = encoded_control[ 14];
   assign decoded_control[ 15] = encoded_control[ 15];
   assign decoded_control[ 16] = encoded_control[ 16];
   assign decoded_control[ 17] = encoded_control[ 17];
   assign decoded_control[ 18] = encoded_control[ 18];
   assign decoded_control[ 19] = encoded_control[ 19];
   assign decoded_control[ 20] = encoded_control[ 20];
   assign decoded_control[ 21] = encoded_control[ 21];
   assign decoded_control[ 22] = encoded_control[ 22];
   assign decoded_control[ 23] = encoded_control[ 23];
   assign decoded_control[ 24] = encoded_control[ 24];
   assign decoded_control[ 25] = encoded_control[ 25];
   assign decoded_control[ 26] = encoded_control[ 26];
   assign decoded_control[ 27] = encoded_control[ 27];
   assign decoded_control[ 28] = encoded_control[ 28];
   assign decoded_control[ 29] = encoded_control[ 29];
   assign decoded_control[ 30] = encoded_control[ 30];
   assign decoded_control[ 31] = encoded_control[ 31];
   assign decoded_control[ 32] = encoded_control[ 32];
   assign decoded_control[ 33] = encoded_control[ 33];
   assign decoded_control[ 34] = encoded_control[ 34];
   assign decoded_control[ 35] = encoded_control[ 35];
   assign decoded_control[ 36] = encoded_control[ 36];
   assign decoded_control[ 37] = encoded_control[ 37];
   assign decoded_control[ 38] = encoded_control[ 38];
   assign decoded_control[ 39] = encoded_control[ 39];
   assign decoded_control[ 40] = encoded_control[ 40];
   assign decoded_control[ 41] = encoded_control[ 41];
   assign decoded_control[ 42] = encoded_control[ 42];
   assign decoded_control[ 43] = encoded_control[ 43];
   assign decoded_control[ 44] = encoded_control[ 44];
   assign decoded_control[ 45] = encoded_control[ 45];
   assign decoded_control[ 46] = encoded_control[ 46];
   assign decoded_control[ 47] = encoded_control[ 47];
   assign decoded_control[ 48] = encoded_control[ 48];
   assign decoded_control[ 49] = encoded_control[ 49];
   assign decoded_control[ 50] = encoded_control[ 50];
   assign decoded_control[ 51] = encoded_control[ 51];
   assign decoded_control[ 52] = encoded_control[ 52];
   assign decoded_control[ 53] = encoded_control[ 53];
   assign decoded_control[ 54] = encoded_control[ 54];
   assign decoded_control[ 55] = encoded_control[ 55];
   assign decoded_control[ 56] = encoded_control[ 56];
   assign decoded_control[ 57] = encoded_control[ 57];
   assign decoded_control[ 58] = encoded_control[ 58];
   assign decoded_control[ 59] = encoded_control[ 59];
   assign decoded_control[ 60] = encoded_control[ 60];
   assign decoded_control[ 61] = encoded_control[ 61];
   assign decoded_control[ 62] = encoded_control[ 62];
   assign decoded_control[ 63] = encoded_control[ 63];
   assign decoded_control[ 64] = encoded_control[ 64];
   assign decoded_control[ 65] = encoded_control[ 65];
   assign decoded_control[ 66] = encoded_control[ 66];
   assign decoded_control[ 67] = encoded_control[ 67];
   assign decoded_control[ 68] = encoded_control[ 68];
   assign decoded_control[ 69] = encoded_control[ 69];
   assign decoded_control[ 70] = encoded_control[ 70];
   assign decoded_control[ 71] = encoded_control[ 71];
   assign decoded_control[ 72] = encoded_control[ 72];
   assign decoded_control[ 73] = encoded_control[ 73];
   assign decoded_control[ 74] = encoded_control[ 74];
   assign decoded_control[ 75] = encoded_control[ 75];
   assign decoded_control[ 76] = encoded_control[ 76];
   assign decoded_control[ 77] = encoded_control[ 77];
   assign decoded_control[ 78] = encoded_control[ 78];
   assign decoded_control[ 79] = encoded_control[ 79];
   assign decoded_control[ 80] = encoded_control[ 80];
   assign decoded_control[ 81] = encoded_control[ 81];
   assign decoded_control[ 82] = encoded_control[ 82];
   assign decoded_control[ 83] = encoded_control[ 83];
   assign decoded_control[ 84] = encoded_control[ 84];
   assign decoded_control[ 85] = encoded_control[ 85];
   assign decoded_control[ 86] = encoded_control[ 86];
   assign decoded_control[ 87] = encoded_control[ 87];
   assign decoded_control[ 88] = encoded_control[ 88];
   assign decoded_control[ 89] = encoded_control[ 89];
   assign decoded_control[ 90] = encoded_control[ 90];
   assign decoded_control[ 91] = encoded_control[ 91];
   assign decoded_control[ 92] = encoded_control[ 92];
   assign decoded_control[ 93] = encoded_control[ 93];
   assign decoded_control[ 94] = encoded_control[ 94];
   assign decoded_control[ 95] = encoded_control[ 95];
   assign decoded_control[ 96] = encoded_control[ 96];
   assign decoded_control[ 97] = encoded_control[ 97];
   assign decoded_control[ 98] = encoded_control[ 98];
   assign decoded_control[ 99] = encoded_control[ 99];
   assign decoded_control[100] = encoded_control[100];
   assign decoded_control[101] = encoded_control[101];
   assign decoded_control[102] = encoded_control[102];
   assign decoded_control[103] = encoded_control[103];
   assign decoded_control[104] = encoded_control[104];
   assign decoded_control[105] = encoded_control[105];
   assign decoded_control[106] = encoded_control[106];
   assign decoded_control[107] = encoded_control[107];
   assign decoded_control[108] = encoded_control[108];
   assign decoded_control[109] = encoded_control[109];
   assign decoded_control[110] = encoded_control[110];
   assign decoded_control[111] = encoded_control[111];
   assign decoded_control[112] = encoded_control[112];
   assign decoded_control[113] = encoded_control[113];
   assign decoded_control[114] = encoded_control[114];
   assign decoded_control[115] = encoded_control[115];
   assign decoded_control[116] = encoded_control[116];
   assign decoded_control[117] = encoded_control[117];
   assign decoded_control[118] = encoded_control[118];
   assign decoded_control[119] = encoded_control[119];
   assign decoded_control[120] = encoded_control[120];
   assign decoded_control[121] = encoded_control[121];
   assign decoded_control[122] = encoded_control[122];
   assign decoded_control[123] = encoded_control[123];
   assign decoded_control[124] = encoded_control[124];
   assign decoded_control[125] = encoded_control[125];
   assign decoded_control[126] = encoded_control[126];
   assign decoded_control[127] = encoded_control[127];
   assign decoded_control[128] = encoded_control[128];
   assign decoded_control[129] = encoded_control[129];
   assign decoded_control[130] = encoded_control[130];
   assign decoded_control[131] = encoded_control[131];
   assign decoded_control[132] = encoded_control[132];
   assign decoded_control[133] = encoded_control[133];
   assign decoded_control[134] = encoded_control[134];
   assign decoded_control[135] = encoded_control[135];
   assign decoded_control[136] = encoded_control[136];
   assign decoded_control[137] = encoded_control[137];
   assign decoded_control[138] = encoded_control[138];
   assign decoded_control[139] = encoded_control[139];
   assign decoded_control[140] = encoded_control[140];
   assign decoded_control[141] = encoded_control[141];
   assign decoded_control[142] = encoded_control[142];
   assign decoded_control[143] = encoded_control[143];
   assign decoded_control[144] = encoded_control[144];
   assign decoded_control[145] = encoded_control[145];
   assign decoded_control[146] = encoded_control[146];
   assign decoded_control[147] = encoded_control[147];
   assign decoded_control[148] = encoded_control[148];
   assign decoded_control[149] = encoded_control[149];
   assign decoded_control[150] = encoded_control[150];
   assign decoded_control[151] = encoded_control[151];
   assign decoded_control[152] = encoded_control[152];
   assign decoded_control[153] = encoded_control[153];
   assign decoded_control[154] = encoded_control[154];
   assign decoded_control[155] = encoded_control[155];
   assign decoded_control[156] = encoded_control[156];
   assign decoded_control[157] = encoded_control[157];
   assign decoded_control[158] = encoded_control[158];
   assign decoded_control[159] = encoded_control[159];
   assign decoded_control[160] = encoded_control[160];
   assign decoded_control[161] = encoded_control[161];
   assign decoded_control[162] = encoded_control[162];
   assign decoded_control[163] = encoded_control[163];
   assign decoded_control[164] = encoded_control[164];
   assign decoded_control[165] = encoded_control[165];
   assign decoded_control[166] = encoded_control[166];
   assign decoded_control[167] = encoded_control[167];
   assign decoded_control[168] = encoded_control[168];
   assign decoded_control[169] = encoded_control[169];
   assign decoded_control[170] = encoded_control[170];
   assign decoded_control[171] = encoded_control[171];
   assign decoded_control[172] = encoded_control[172];
   assign decoded_control[173] = encoded_control[173];
   assign decoded_control[174] = encoded_control[174];
   assign decoded_control[175] = encoded_control[175];
   assign decoded_control[176] = encoded_control[176];
   assign decoded_control[177] = encoded_control[177];
   assign decoded_control[178] = encoded_control[178];
   assign decoded_control[179] = encoded_control[179];
   assign decoded_control[180] = encoded_control[180];
   assign decoded_control[181] = encoded_control[181];
   assign decoded_control[182] = encoded_control[182];
   assign decoded_control[183] = encoded_control[183];
   assign decoded_control[184] = encoded_control[184];
   assign decoded_control[185] = encoded_control[185];
   assign decoded_control[186] = encoded_control[186];
   assign decoded_control[187] = encoded_control[187];
   assign decoded_control[188] = encoded_control[188];
   assign decoded_control[189] = encoded_control[189];
   assign decoded_control[190] = encoded_control[190];
   assign decoded_control[191] = encoded_control[191];
   assign decoded_control[192] = encoded_control[192];
   assign decoded_control[193] = encoded_control[193];
   assign decoded_control[194] = encoded_control[194];
   assign decoded_control[195] = encoded_control[195];
   assign decoded_control[196] = encoded_control[196];
   assign decoded_control[197] = encoded_control[197];
   assign decoded_control[198] = encoded_control[198];
   assign decoded_control[199] = encoded_control[199];
   assign decoded_control[200] = encoded_control[200];
   assign decoded_control[201] = encoded_control[201];
   assign decoded_control[202] = encoded_control[202];
   assign decoded_control[203] = encoded_control[203];
   assign decoded_control[204] = encoded_control[204];
   assign decoded_control[205] = encoded_control[205];
   assign decoded_control[206] = encoded_control[206];
   assign decoded_control[207] = encoded_control[207];
   assign decoded_control[208] = encoded_control[208];
   assign decoded_control[209] = encoded_control[209];
   assign decoded_control[210] = encoded_control[210];
   assign decoded_control[211] = encoded_control[211];
   assign decoded_control[212] = encoded_control[212];
   assign decoded_control[213] = encoded_control[213];
   assign decoded_control[214] = encoded_control[214];
   assign decoded_control[215] = encoded_control[215];
   assign decoded_control[216] = encoded_control[216];
   assign decoded_control[217] = encoded_control[217];
   assign decoded_control[218] = encoded_control[218];
   assign decoded_control[219] = encoded_control[219];
   assign decoded_control[220] = encoded_control[220];
   assign decoded_control[221] = encoded_control[221];
   assign decoded_control[222] = encoded_control[222];
   assign decoded_control[223] = encoded_control[223];
   assign decoded_control[224] = encoded_control[224];
   assign decoded_control[225] = encoded_control[225];
   assign decoded_control[226] = encoded_control[226];
   assign decoded_control[227] = encoded_control[227];
   assign decoded_control[228] = encoded_control[228];
   assign decoded_control[229] = encoded_control[229];
   assign decoded_control[230] = encoded_control[230];
   assign decoded_control[231] = encoded_control[231];
   assign decoded_control[232] = encoded_control[232];
   assign decoded_control[233] = encoded_control[233];
   assign decoded_control[234] = encoded_control[234];
   assign decoded_control[235] = encoded_control[235];
   assign decoded_control[236] = encoded_control[236];
   assign decoded_control[237] = encoded_control[237];
   assign decoded_control[238] = encoded_control[238];
   assign decoded_control[239] = encoded_control[239];
   assign decoded_control[240] = encoded_control[240];
   assign decoded_control[241] = encoded_control[241];
   assign decoded_control[242] = encoded_control[242];
   assign decoded_control[243] = encoded_control[243];
   assign decoded_control[244] = encoded_control[244];
   assign decoded_control[245] = encoded_control[245];
   assign decoded_control[246] = encoded_control[246];
   assign decoded_control[247] = encoded_control[247];
   assign decoded_control[248] = encoded_control[248];
   assign decoded_control[249] = encoded_control[249];
   assign decoded_control[250] = encoded_control[250];
   assign decoded_control[251] = encoded_control[251];
   assign decoded_control[252] = encoded_control[252];
   assign decoded_control[253] = encoded_control[253];
   assign decoded_control[254] = encoded_control[254];
   assign decoded_control[255] = encoded_control[255];
   assign decoded_control[256] = encoded_control[256];
   assign decoded_control[257] = encoded_control[257];
   assign decoded_control[258] = encoded_control[258];
   assign decoded_control[259] = encoded_control[259];
   assign decoded_control[260] = encoded_control[260];
   assign decoded_control[261] = encoded_control[261];
   assign decoded_control[262] = encoded_control[262];
   assign decoded_control[263] = encoded_control[263];
   assign decoded_control[264] = encoded_control[264];
   assign decoded_control[265] = encoded_control[265];
   assign decoded_control[266] = encoded_control[266];
   assign decoded_control[267] = encoded_control[267];
   assign decoded_control[268] = encoded_control[268];
   assign decoded_control[269] = encoded_control[269];
   assign decoded_control[270] = encoded_control[270];
   assign decoded_control[271] = encoded_control[271];
   assign decoded_control[272] = encoded_control[272];
   assign decoded_control[273] = encoded_control[273];
   assign decoded_control[274] = encoded_control[274];
   assign decoded_control[275] = encoded_control[275];
   assign decoded_control[276] = encoded_control[276];
   assign decoded_control[277] = encoded_control[277];
   assign decoded_control[278] = encoded_control[278];
   assign decoded_control[279] = encoded_control[279];
   assign decoded_control[280] = encoded_control[280];
   assign decoded_control[281] = encoded_control[281];
   assign decoded_control[282] = encoded_control[282];
   assign decoded_control[283] = encoded_control[283];
   assign decoded_control[284] = encoded_control[284];
   assign decoded_control[285] = encoded_control[285];
   assign decoded_control[286] = encoded_control[286];
   assign decoded_control[287] = encoded_control[287];
   assign decoded_control[288] = encoded_control[288];
   assign decoded_control[289] = encoded_control[289];
   assign decoded_control[290] = encoded_control[290];
   assign decoded_control[291] = encoded_control[291];
   assign decoded_control[292] = encoded_control[292];
   assign decoded_control[293] = encoded_control[293];
   assign decoded_control[294] = encoded_control[294];
   assign decoded_control[295] = encoded_control[295];
   assign decoded_control[296] = encoded_control[296];
   assign decoded_control[297] = encoded_control[297];
   assign decoded_control[298] = encoded_control[298];
   assign decoded_control[299] = encoded_control[299];
   assign decoded_control[300] = encoded_control[300];
   assign decoded_control[301] = encoded_control[301];
   assign decoded_control[302] = encoded_control[302];
   assign decoded_control[303] = encoded_control[303];
   assign decoded_control[304] = encoded_control[304];
   assign decoded_control[305] = encoded_control[305];
   assign decoded_control[306] = encoded_control[306];
   assign decoded_control[307] = encoded_control[307];
   assign decoded_control[308] = encoded_control[308];
   assign decoded_control[309] = encoded_control[309];
   assign decoded_control[310] = encoded_control[310];
   assign decoded_control[311] = encoded_control[311];
   assign decoded_control[312] = encoded_control[312];
   assign decoded_control[313] = encoded_control[313];
   assign decoded_control[314] = encoded_control[314];
   assign decoded_control[315] = encoded_control[315];
   assign decoded_control[316] = encoded_control[316];
   assign decoded_control[317] = encoded_control[317];
   assign decoded_control[318] = encoded_control[318];
   assign decoded_control[319] = encoded_control[319];
   assign decoded_control[320] = encoded_control[320];
   assign decoded_control[321] = encoded_control[321];
   assign decoded_control[322] = encoded_control[322];
   assign decoded_control[323] = encoded_control[323];
   assign decoded_control[324] = encoded_control[324];
   assign decoded_control[325] = encoded_control[325];
   assign decoded_control[326] = encoded_control[326];
   assign decoded_control[327] = encoded_control[327];
   assign decoded_control[328] = encoded_control[328];
   assign decoded_control[329] = encoded_control[329];
   assign decoded_control[330] = encoded_control[330];
   assign decoded_control[331] = encoded_control[331];
   assign decoded_control[332] = encoded_control[332];
   assign decoded_control[333] = encoded_control[333];
   assign decoded_control[334] = encoded_control[334];
   assign decoded_control[335] = encoded_control[335];
   assign decoded_control[336] = encoded_control[336];
   assign decoded_control[337] = encoded_control[337];
   assign decoded_control[338] = encoded_control[338];
   assign decoded_control[339] = encoded_control[339];
   assign decoded_control[340] = encoded_control[340];
   assign decoded_control[341] = encoded_control[341];
   assign decoded_control[342] = encoded_control[342];
   assign decoded_control[343] = encoded_control[343];
   assign decoded_control[344] = encoded_control[344];
   assign decoded_control[345] = encoded_control[345];
   assign decoded_control[346] = encoded_control[346];
   assign decoded_control[347] = encoded_control[347];
   assign decoded_control[348] = encoded_control[348];
   assign decoded_control[349] = encoded_control[349];
   assign decoded_control[350] = encoded_control[350];
   assign decoded_control[351] = encoded_control[351];
   assign decoded_control[352] = encoded_control[352];
   assign decoded_control[353] = encoded_control[353];
   assign decoded_control[354] = encoded_control[354];
   assign decoded_control[355] = encoded_control[355];
   assign decoded_control[356] = encoded_control[356];
   assign decoded_control[357] = encoded_control[357];
   assign decoded_control[358] = encoded_control[358];
   assign decoded_control[359] = encoded_control[359];
   assign decoded_control[360] = encoded_control[360];
   assign decoded_control[361] = encoded_control[361];
   assign decoded_control[362] = encoded_control[362];
   assign decoded_control[363] = encoded_control[363];
   assign decoded_control[364] = encoded_control[364];
   assign decoded_control[365] = encoded_control[365];
   assign decoded_control[366] = encoded_control[366];
   assign decoded_control[367] = encoded_control[367];
   assign decoded_control[368] = encoded_control[368];
   assign decoded_control[369] = encoded_control[369];
   assign decoded_control[370] = encoded_control[370];
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_low_power_shift_controller (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire         edt_low_power_shift_en,
   input  wire [  3:0] edt_channels_in,
   input  wire [370:0] edt_decompressor_out,
   output wire [  3:0] edt_channels_out_from_low_power_shift_control,
   output wire [370:0] edt_scan_in
);
   reg    [ 92:0] low_power_shift_reg_0;
   reg    [ 92:0] low_power_shift_reg_1;
   reg    [ 92:0] low_power_shift_reg_2;
   reg    [ 91:0] low_power_shift_reg_3;
   reg    [ 92:0] low_power_hold_reg_0;
   reg    [ 92:0] low_power_hold_reg_1;
   reg    [ 92:0] low_power_hold_reg_2;
   reg    [ 91:0] low_power_hold_reg_3;
   wire   [370:0] encoded_control;
   wire   [370:0] bias_inputs;
   wire           low_power_shift_reg_sync_reset;
   wire           low_power_hold_reg_sync_set;

   assign low_power_shift_reg_sync_reset = edt_update;

   // synopsys sync_set_reset low_power_shift_reg_sync_reset
   always @(posedge edt_clock)
   begin : shift_low_power_regs
      if (low_power_shift_reg_sync_reset == 1'b1) begin
         low_power_shift_reg_0 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         low_power_shift_reg_1 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         low_power_shift_reg_2 <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         low_power_shift_reg_3 <= 92'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      end
      else begin
         low_power_shift_reg_0 <= {edt_channels_in[0], low_power_shift_reg_0[92:1]};
         low_power_shift_reg_1 <= {edt_channels_in[1], low_power_shift_reg_1[92:1]};
         low_power_shift_reg_2 <= {edt_channels_in[2], low_power_shift_reg_2[92:1]};
         low_power_shift_reg_3 <= {edt_channels_in[3], low_power_shift_reg_3[91:1]};
      end
   end

   assign low_power_hold_reg_sync_set = edt_update & ~edt_low_power_shift_en;

   // synopsys sync_set_reset low_power_hold_reg_sync_set
   always @(posedge edt_clock)
   begin : update_low_power_regs
      if (low_power_hold_reg_sync_set == 1'b1) begin
         low_power_hold_reg_0 <= 93'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
         low_power_hold_reg_1 <= 93'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
         low_power_hold_reg_2 <= 93'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
         low_power_hold_reg_3 <= 92'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
      end
      else begin
         if (edt_update == 1'b1) begin
            low_power_hold_reg_0 <= low_power_shift_reg_0;
            low_power_hold_reg_1 <= low_power_shift_reg_1;
            low_power_hold_reg_2 <= low_power_shift_reg_2;
            low_power_hold_reg_3 <= low_power_shift_reg_3;
         end
      end
   end

   assign edt_channels_out_from_low_power_shift_control[0] = edt_low_power_shift_en ? low_power_shift_reg_0[0] : edt_channels_in[0];
   assign edt_channels_out_from_low_power_shift_control[1] = edt_low_power_shift_en ? low_power_shift_reg_1[0] : edt_channels_in[1];
   assign edt_channels_out_from_low_power_shift_control[2] = edt_low_power_shift_en ? low_power_shift_reg_2[0] : edt_channels_in[2];
   assign edt_channels_out_from_low_power_shift_control[3] = edt_low_power_shift_en ? low_power_shift_reg_3[0] : edt_channels_in[3];

   assign encoded_control = {low_power_hold_reg_3[91], low_power_hold_reg_3[90], low_power_hold_reg_3[89], 
                             low_power_hold_reg_3[88], low_power_hold_reg_3[87], low_power_hold_reg_3[86], 
                             low_power_hold_reg_3[85], low_power_hold_reg_3[84], low_power_hold_reg_3[83], 
                             low_power_hold_reg_3[82], low_power_hold_reg_3[81], low_power_hold_reg_3[80], 
                             low_power_hold_reg_3[79], low_power_hold_reg_3[78], low_power_hold_reg_3[77], 
                             low_power_hold_reg_3[76], low_power_hold_reg_3[75], low_power_hold_reg_3[74], 
                             low_power_hold_reg_3[73], low_power_hold_reg_3[72], low_power_hold_reg_3[71], 
                             low_power_hold_reg_3[70], low_power_hold_reg_3[69], low_power_hold_reg_3[68], 
                             low_power_hold_reg_3[67], low_power_hold_reg_3[66], low_power_hold_reg_3[65], 
                             low_power_hold_reg_3[64], low_power_hold_reg_3[63], low_power_hold_reg_3[62], 
                             low_power_hold_reg_3[61], low_power_hold_reg_3[60], low_power_hold_reg_3[59], 
                             low_power_hold_reg_3[58], low_power_hold_reg_3[57], low_power_hold_reg_3[56], 
                             low_power_hold_reg_3[55], low_power_hold_reg_3[54], low_power_hold_reg_3[53], 
                             low_power_hold_reg_3[52], low_power_hold_reg_3[51], low_power_hold_reg_3[50], 
                             low_power_hold_reg_3[49], low_power_hold_reg_3[48], low_power_hold_reg_3[47], 
                             low_power_hold_reg_3[46], low_power_hold_reg_3[45], low_power_hold_reg_3[44], 
                             low_power_hold_reg_3[43], low_power_hold_reg_3[42], low_power_hold_reg_3[41], 
                             low_power_hold_reg_3[40], low_power_hold_reg_3[39], low_power_hold_reg_3[38], 
                             low_power_hold_reg_3[37], low_power_hold_reg_3[36], low_power_hold_reg_3[35], 
                             low_power_hold_reg_3[34], low_power_hold_reg_3[33], low_power_hold_reg_3[32], 
                             low_power_hold_reg_3[31], low_power_hold_reg_3[30], low_power_hold_reg_3[29], 
                             low_power_hold_reg_3[28], low_power_hold_reg_3[27], low_power_hold_reg_3[26], 
                             low_power_hold_reg_3[25], low_power_hold_reg_3[24], low_power_hold_reg_3[23], 
                             low_power_hold_reg_3[22], low_power_hold_reg_3[21], low_power_hold_reg_3[20], 
                             low_power_hold_reg_3[19], low_power_hold_reg_3[18], low_power_hold_reg_3[17], 
                             low_power_hold_reg_3[16], low_power_hold_reg_3[15], low_power_hold_reg_3[14], 
                             low_power_hold_reg_3[13], low_power_hold_reg_3[12], low_power_hold_reg_3[11], 
                             low_power_hold_reg_3[10], low_power_hold_reg_3[9], low_power_hold_reg_3[8], 
                             low_power_hold_reg_3[7], low_power_hold_reg_3[6], low_power_hold_reg_3[5], 
                             low_power_hold_reg_3[4], low_power_hold_reg_3[3], low_power_hold_reg_3[2], 
                             low_power_hold_reg_3[1], low_power_hold_reg_3[0], low_power_hold_reg_2[92], 
                             low_power_hold_reg_2[91], low_power_hold_reg_2[90], low_power_hold_reg_2[89], 
                             low_power_hold_reg_2[88], low_power_hold_reg_2[87], low_power_hold_reg_2[86], 
                             low_power_hold_reg_2[85], low_power_hold_reg_2[84], low_power_hold_reg_2[83], 
                             low_power_hold_reg_2[82], low_power_hold_reg_2[81], low_power_hold_reg_2[80], 
                             low_power_hold_reg_2[79], low_power_hold_reg_2[78], low_power_hold_reg_2[77], 
                             low_power_hold_reg_2[76], low_power_hold_reg_2[75], low_power_hold_reg_2[74], 
                             low_power_hold_reg_2[73], low_power_hold_reg_2[72], low_power_hold_reg_2[71], 
                             low_power_hold_reg_2[70], low_power_hold_reg_2[69], low_power_hold_reg_2[68], 
                             low_power_hold_reg_2[67], low_power_hold_reg_2[66], low_power_hold_reg_2[65], 
                             low_power_hold_reg_2[64], low_power_hold_reg_2[63], low_power_hold_reg_2[62], 
                             low_power_hold_reg_2[61], low_power_hold_reg_2[60], low_power_hold_reg_2[59], 
                             low_power_hold_reg_2[58], low_power_hold_reg_2[57], low_power_hold_reg_2[56], 
                             low_power_hold_reg_2[55], low_power_hold_reg_2[54], low_power_hold_reg_2[53], 
                             low_power_hold_reg_2[52], low_power_hold_reg_2[51], low_power_hold_reg_2[50], 
                             low_power_hold_reg_2[49], low_power_hold_reg_2[48], low_power_hold_reg_2[47], 
                             low_power_hold_reg_2[46], low_power_hold_reg_2[45], low_power_hold_reg_2[44], 
                             low_power_hold_reg_2[43], low_power_hold_reg_2[42], low_power_hold_reg_2[41], 
                             low_power_hold_reg_2[40], low_power_hold_reg_2[39], low_power_hold_reg_2[38], 
                             low_power_hold_reg_2[37], low_power_hold_reg_2[36], low_power_hold_reg_2[35], 
                             low_power_hold_reg_2[34], low_power_hold_reg_2[33], low_power_hold_reg_2[32], 
                             low_power_hold_reg_2[31], low_power_hold_reg_2[30], low_power_hold_reg_2[29], 
                             low_power_hold_reg_2[28], low_power_hold_reg_2[27], low_power_hold_reg_2[26], 
                             low_power_hold_reg_2[25], low_power_hold_reg_2[24], low_power_hold_reg_2[23], 
                             low_power_hold_reg_2[22], low_power_hold_reg_2[21], low_power_hold_reg_2[20], 
                             low_power_hold_reg_2[19], low_power_hold_reg_2[18], low_power_hold_reg_2[17], 
                             low_power_hold_reg_2[16], low_power_hold_reg_2[15], low_power_hold_reg_2[14], 
                             low_power_hold_reg_2[13], low_power_hold_reg_2[12], low_power_hold_reg_2[11], 
                             low_power_hold_reg_2[10], low_power_hold_reg_2[9], low_power_hold_reg_2[8], 
                             low_power_hold_reg_2[7], low_power_hold_reg_2[6], low_power_hold_reg_2[5], 
                             low_power_hold_reg_2[4], low_power_hold_reg_2[3], low_power_hold_reg_2[2], 
                             low_power_hold_reg_2[1], low_power_hold_reg_2[0], low_power_hold_reg_1[92], 
                             low_power_hold_reg_1[91], low_power_hold_reg_1[90], low_power_hold_reg_1[89], 
                             low_power_hold_reg_1[88], low_power_hold_reg_1[87], low_power_hold_reg_1[86], 
                             low_power_hold_reg_1[85], low_power_hold_reg_1[84], low_power_hold_reg_1[83], 
                             low_power_hold_reg_1[82], low_power_hold_reg_1[81], low_power_hold_reg_1[80], 
                             low_power_hold_reg_1[79], low_power_hold_reg_1[78], low_power_hold_reg_1[77], 
                             low_power_hold_reg_1[76], low_power_hold_reg_1[75], low_power_hold_reg_1[74], 
                             low_power_hold_reg_1[73], low_power_hold_reg_1[72], low_power_hold_reg_1[71], 
                             low_power_hold_reg_1[70], low_power_hold_reg_1[69], low_power_hold_reg_1[68], 
                             low_power_hold_reg_1[67], low_power_hold_reg_1[66], low_power_hold_reg_1[65], 
                             low_power_hold_reg_1[64], low_power_hold_reg_1[63], low_power_hold_reg_1[62], 
                             low_power_hold_reg_1[61], low_power_hold_reg_1[60], low_power_hold_reg_1[59], 
                             low_power_hold_reg_1[58], low_power_hold_reg_1[57], low_power_hold_reg_1[56], 
                             low_power_hold_reg_1[55], low_power_hold_reg_1[54], low_power_hold_reg_1[53], 
                             low_power_hold_reg_1[52], low_power_hold_reg_1[51], low_power_hold_reg_1[50], 
                             low_power_hold_reg_1[49], low_power_hold_reg_1[48], low_power_hold_reg_1[47], 
                             low_power_hold_reg_1[46], low_power_hold_reg_1[45], low_power_hold_reg_1[44], 
                             low_power_hold_reg_1[43], low_power_hold_reg_1[42], low_power_hold_reg_1[41], 
                             low_power_hold_reg_1[40], low_power_hold_reg_1[39], low_power_hold_reg_1[38], 
                             low_power_hold_reg_1[37], low_power_hold_reg_1[36], low_power_hold_reg_1[35], 
                             low_power_hold_reg_1[34], low_power_hold_reg_1[33], low_power_hold_reg_1[32], 
                             low_power_hold_reg_1[31], low_power_hold_reg_1[30], low_power_hold_reg_1[29], 
                             low_power_hold_reg_1[28], low_power_hold_reg_1[27], low_power_hold_reg_1[26], 
                             low_power_hold_reg_1[25], low_power_hold_reg_1[24], low_power_hold_reg_1[23], 
                             low_power_hold_reg_1[22], low_power_hold_reg_1[21], low_power_hold_reg_1[20], 
                             low_power_hold_reg_1[19], low_power_hold_reg_1[18], low_power_hold_reg_1[17], 
                             low_power_hold_reg_1[16], low_power_hold_reg_1[15], low_power_hold_reg_1[14], 
                             low_power_hold_reg_1[13], low_power_hold_reg_1[12], low_power_hold_reg_1[11], 
                             low_power_hold_reg_1[10], low_power_hold_reg_1[9], low_power_hold_reg_1[8], 
                             low_power_hold_reg_1[7], low_power_hold_reg_1[6], low_power_hold_reg_1[5], 
                             low_power_hold_reg_1[4], low_power_hold_reg_1[3], low_power_hold_reg_1[2], 
                             low_power_hold_reg_1[1], low_power_hold_reg_1[0], low_power_hold_reg_0[92], 
                             low_power_hold_reg_0[91], low_power_hold_reg_0[90], low_power_hold_reg_0[89], 
                             low_power_hold_reg_0[88], low_power_hold_reg_0[87], low_power_hold_reg_0[86], 
                             low_power_hold_reg_0[85], low_power_hold_reg_0[84], low_power_hold_reg_0[83], 
                             low_power_hold_reg_0[82], low_power_hold_reg_0[81], low_power_hold_reg_0[80], 
                             low_power_hold_reg_0[79], low_power_hold_reg_0[78], low_power_hold_reg_0[77], 
                             low_power_hold_reg_0[76], low_power_hold_reg_0[75], low_power_hold_reg_0[74], 
                             low_power_hold_reg_0[73], low_power_hold_reg_0[72], low_power_hold_reg_0[71], 
                             low_power_hold_reg_0[70], low_power_hold_reg_0[69], low_power_hold_reg_0[68], 
                             low_power_hold_reg_0[67], low_power_hold_reg_0[66], low_power_hold_reg_0[65], 
                             low_power_hold_reg_0[64], low_power_hold_reg_0[63], low_power_hold_reg_0[62], 
                             low_power_hold_reg_0[61], low_power_hold_reg_0[60], low_power_hold_reg_0[59], 
                             low_power_hold_reg_0[58], low_power_hold_reg_0[57], low_power_hold_reg_0[56], 
                             low_power_hold_reg_0[55], low_power_hold_reg_0[54], low_power_hold_reg_0[53], 
                             low_power_hold_reg_0[52], low_power_hold_reg_0[51], low_power_hold_reg_0[50], 
                             low_power_hold_reg_0[49], low_power_hold_reg_0[48], low_power_hold_reg_0[47], 
                             low_power_hold_reg_0[46], low_power_hold_reg_0[45], low_power_hold_reg_0[44], 
                             low_power_hold_reg_0[43], low_power_hold_reg_0[42], low_power_hold_reg_0[41], 
                             low_power_hold_reg_0[40], low_power_hold_reg_0[39], low_power_hold_reg_0[38], 
                             low_power_hold_reg_0[37], low_power_hold_reg_0[36], low_power_hold_reg_0[35], 
                             low_power_hold_reg_0[34], low_power_hold_reg_0[33], low_power_hold_reg_0[32], 
                             low_power_hold_reg_0[31], low_power_hold_reg_0[30], low_power_hold_reg_0[29], 
                             low_power_hold_reg_0[28], low_power_hold_reg_0[27], low_power_hold_reg_0[26], 
                             low_power_hold_reg_0[25], low_power_hold_reg_0[24], low_power_hold_reg_0[23], 
                             low_power_hold_reg_0[22], low_power_hold_reg_0[21], low_power_hold_reg_0[20], 
                             low_power_hold_reg_0[19], low_power_hold_reg_0[18], low_power_hold_reg_0[17], 
                             low_power_hold_reg_0[16], low_power_hold_reg_0[15], low_power_hold_reg_0[14], 
                             low_power_hold_reg_0[13], low_power_hold_reg_0[12], low_power_hold_reg_0[11], 
                             low_power_hold_reg_0[10], low_power_hold_reg_0[9], low_power_hold_reg_0[8], 
                             low_power_hold_reg_0[7], low_power_hold_reg_0[6], low_power_hold_reg_0[5], 
                             low_power_hold_reg_0[4], low_power_hold_reg_0[3], low_power_hold_reg_0[2], 
                             low_power_hold_reg_0[1], low_power_hold_reg_0[0]};

   firebird7_in_gate2_tessent_edt_intest_edt_low_power_shift_decoder decoder (
      .encoded_control(encoded_control),
      .decoded_control(bias_inputs));

   assign edt_scan_in[  0] = edt_decompressor_out[  0] & bias_inputs[  0];
   assign edt_scan_in[  1] = edt_decompressor_out[  1] & bias_inputs[  1];
   assign edt_scan_in[  2] = edt_decompressor_out[  2] & bias_inputs[  2];
   assign edt_scan_in[  3] = edt_decompressor_out[  3] & bias_inputs[  3];
   assign edt_scan_in[  4] = edt_decompressor_out[  4] & bias_inputs[  4];
   assign edt_scan_in[  5] = edt_decompressor_out[  5] & bias_inputs[  5];
   assign edt_scan_in[  6] = edt_decompressor_out[  6] & bias_inputs[  6];
   assign edt_scan_in[  7] = edt_decompressor_out[  7] & bias_inputs[  7];
   assign edt_scan_in[  8] = edt_decompressor_out[  8] & bias_inputs[  8];
   assign edt_scan_in[  9] = edt_decompressor_out[  9] & bias_inputs[  9];
   assign edt_scan_in[ 10] = edt_decompressor_out[ 10] & bias_inputs[ 10];
   assign edt_scan_in[ 11] = edt_decompressor_out[ 11] & bias_inputs[ 11];
   assign edt_scan_in[ 12] = edt_decompressor_out[ 12] & bias_inputs[ 12];
   assign edt_scan_in[ 13] = edt_decompressor_out[ 13] & bias_inputs[ 13];
   assign edt_scan_in[ 14] = edt_decompressor_out[ 14] & bias_inputs[ 14];
   assign edt_scan_in[ 15] = edt_decompressor_out[ 15] & bias_inputs[ 15];
   assign edt_scan_in[ 16] = edt_decompressor_out[ 16] & bias_inputs[ 16];
   assign edt_scan_in[ 17] = edt_decompressor_out[ 17] & bias_inputs[ 17];
   assign edt_scan_in[ 18] = edt_decompressor_out[ 18] & bias_inputs[ 18];
   assign edt_scan_in[ 19] = edt_decompressor_out[ 19] & bias_inputs[ 19];
   assign edt_scan_in[ 20] = edt_decompressor_out[ 20] & bias_inputs[ 20];
   assign edt_scan_in[ 21] = edt_decompressor_out[ 21] & bias_inputs[ 21];
   assign edt_scan_in[ 22] = edt_decompressor_out[ 22] & bias_inputs[ 22];
   assign edt_scan_in[ 23] = edt_decompressor_out[ 23] & bias_inputs[ 23];
   assign edt_scan_in[ 24] = edt_decompressor_out[ 24] & bias_inputs[ 24];
   assign edt_scan_in[ 25] = edt_decompressor_out[ 25] & bias_inputs[ 25];
   assign edt_scan_in[ 26] = edt_decompressor_out[ 26] & bias_inputs[ 26];
   assign edt_scan_in[ 27] = edt_decompressor_out[ 27] & bias_inputs[ 27];
   assign edt_scan_in[ 28] = edt_decompressor_out[ 28] & bias_inputs[ 28];
   assign edt_scan_in[ 29] = edt_decompressor_out[ 29] & bias_inputs[ 29];
   assign edt_scan_in[ 30] = edt_decompressor_out[ 30] & bias_inputs[ 30];
   assign edt_scan_in[ 31] = edt_decompressor_out[ 31] & bias_inputs[ 31];
   assign edt_scan_in[ 32] = edt_decompressor_out[ 32] & bias_inputs[ 32];
   assign edt_scan_in[ 33] = edt_decompressor_out[ 33] & bias_inputs[ 33];
   assign edt_scan_in[ 34] = edt_decompressor_out[ 34] & bias_inputs[ 34];
   assign edt_scan_in[ 35] = edt_decompressor_out[ 35] & bias_inputs[ 35];
   assign edt_scan_in[ 36] = edt_decompressor_out[ 36] & bias_inputs[ 36];
   assign edt_scan_in[ 37] = edt_decompressor_out[ 37] & bias_inputs[ 37];
   assign edt_scan_in[ 38] = edt_decompressor_out[ 38] & bias_inputs[ 38];
   assign edt_scan_in[ 39] = edt_decompressor_out[ 39] & bias_inputs[ 39];
   assign edt_scan_in[ 40] = edt_decompressor_out[ 40] & bias_inputs[ 40];
   assign edt_scan_in[ 41] = edt_decompressor_out[ 41] & bias_inputs[ 41];
   assign edt_scan_in[ 42] = edt_decompressor_out[ 42] & bias_inputs[ 42];
   assign edt_scan_in[ 43] = edt_decompressor_out[ 43] & bias_inputs[ 43];
   assign edt_scan_in[ 44] = edt_decompressor_out[ 44] & bias_inputs[ 44];
   assign edt_scan_in[ 45] = edt_decompressor_out[ 45] & bias_inputs[ 45];
   assign edt_scan_in[ 46] = edt_decompressor_out[ 46] & bias_inputs[ 46];
   assign edt_scan_in[ 47] = edt_decompressor_out[ 47] & bias_inputs[ 47];
   assign edt_scan_in[ 48] = edt_decompressor_out[ 48] & bias_inputs[ 48];
   assign edt_scan_in[ 49] = edt_decompressor_out[ 49] & bias_inputs[ 49];
   assign edt_scan_in[ 50] = edt_decompressor_out[ 50] & bias_inputs[ 50];
   assign edt_scan_in[ 51] = edt_decompressor_out[ 51] & bias_inputs[ 51];
   assign edt_scan_in[ 52] = edt_decompressor_out[ 52] & bias_inputs[ 52];
   assign edt_scan_in[ 53] = edt_decompressor_out[ 53] & bias_inputs[ 53];
   assign edt_scan_in[ 54] = edt_decompressor_out[ 54] & bias_inputs[ 54];
   assign edt_scan_in[ 55] = edt_decompressor_out[ 55] & bias_inputs[ 55];
   assign edt_scan_in[ 56] = edt_decompressor_out[ 56] & bias_inputs[ 56];
   assign edt_scan_in[ 57] = edt_decompressor_out[ 57] & bias_inputs[ 57];
   assign edt_scan_in[ 58] = edt_decompressor_out[ 58] & bias_inputs[ 58];
   assign edt_scan_in[ 59] = edt_decompressor_out[ 59] & bias_inputs[ 59];
   assign edt_scan_in[ 60] = edt_decompressor_out[ 60] & bias_inputs[ 60];
   assign edt_scan_in[ 61] = edt_decompressor_out[ 61] & bias_inputs[ 61];
   assign edt_scan_in[ 62] = edt_decompressor_out[ 62] & bias_inputs[ 62];
   assign edt_scan_in[ 63] = edt_decompressor_out[ 63] & bias_inputs[ 63];
   assign edt_scan_in[ 64] = edt_decompressor_out[ 64] & bias_inputs[ 64];
   assign edt_scan_in[ 65] = edt_decompressor_out[ 65] & bias_inputs[ 65];
   assign edt_scan_in[ 66] = edt_decompressor_out[ 66] & bias_inputs[ 66];
   assign edt_scan_in[ 67] = edt_decompressor_out[ 67] & bias_inputs[ 67];
   assign edt_scan_in[ 68] = edt_decompressor_out[ 68] & bias_inputs[ 68];
   assign edt_scan_in[ 69] = edt_decompressor_out[ 69] & bias_inputs[ 69];
   assign edt_scan_in[ 70] = edt_decompressor_out[ 70] & bias_inputs[ 70];
   assign edt_scan_in[ 71] = edt_decompressor_out[ 71] & bias_inputs[ 71];
   assign edt_scan_in[ 72] = edt_decompressor_out[ 72] & bias_inputs[ 72];
   assign edt_scan_in[ 73] = edt_decompressor_out[ 73] & bias_inputs[ 73];
   assign edt_scan_in[ 74] = edt_decompressor_out[ 74] & bias_inputs[ 74];
   assign edt_scan_in[ 75] = edt_decompressor_out[ 75] & bias_inputs[ 75];
   assign edt_scan_in[ 76] = edt_decompressor_out[ 76] & bias_inputs[ 76];
   assign edt_scan_in[ 77] = edt_decompressor_out[ 77] & bias_inputs[ 77];
   assign edt_scan_in[ 78] = edt_decompressor_out[ 78] & bias_inputs[ 78];
   assign edt_scan_in[ 79] = edt_decompressor_out[ 79] & bias_inputs[ 79];
   assign edt_scan_in[ 80] = edt_decompressor_out[ 80] & bias_inputs[ 80];
   assign edt_scan_in[ 81] = edt_decompressor_out[ 81] & bias_inputs[ 81];
   assign edt_scan_in[ 82] = edt_decompressor_out[ 82] & bias_inputs[ 82];
   assign edt_scan_in[ 83] = edt_decompressor_out[ 83] & bias_inputs[ 83];
   assign edt_scan_in[ 84] = edt_decompressor_out[ 84] & bias_inputs[ 84];
   assign edt_scan_in[ 85] = edt_decompressor_out[ 85] & bias_inputs[ 85];
   assign edt_scan_in[ 86] = edt_decompressor_out[ 86] & bias_inputs[ 86];
   assign edt_scan_in[ 87] = edt_decompressor_out[ 87] & bias_inputs[ 87];
   assign edt_scan_in[ 88] = edt_decompressor_out[ 88] & bias_inputs[ 88];
   assign edt_scan_in[ 89] = edt_decompressor_out[ 89] & bias_inputs[ 89];
   assign edt_scan_in[ 90] = edt_decompressor_out[ 90] & bias_inputs[ 90];
   assign edt_scan_in[ 91] = edt_decompressor_out[ 91] & bias_inputs[ 91];
   assign edt_scan_in[ 92] = edt_decompressor_out[ 92] & bias_inputs[ 92];
   assign edt_scan_in[ 93] = edt_decompressor_out[ 93] & bias_inputs[ 93];
   assign edt_scan_in[ 94] = edt_decompressor_out[ 94] & bias_inputs[ 94];
   assign edt_scan_in[ 95] = edt_decompressor_out[ 95] & bias_inputs[ 95];
   assign edt_scan_in[ 96] = edt_decompressor_out[ 96] & bias_inputs[ 96];
   assign edt_scan_in[ 97] = edt_decompressor_out[ 97] & bias_inputs[ 97];
   assign edt_scan_in[ 98] = edt_decompressor_out[ 98] & bias_inputs[ 98];
   assign edt_scan_in[ 99] = edt_decompressor_out[ 99] & bias_inputs[ 99];
   assign edt_scan_in[100] = edt_decompressor_out[100] & bias_inputs[100];
   assign edt_scan_in[101] = edt_decompressor_out[101] & bias_inputs[101];
   assign edt_scan_in[102] = edt_decompressor_out[102] & bias_inputs[102];
   assign edt_scan_in[103] = edt_decompressor_out[103] & bias_inputs[103];
   assign edt_scan_in[104] = edt_decompressor_out[104] & bias_inputs[104];
   assign edt_scan_in[105] = edt_decompressor_out[105] & bias_inputs[105];
   assign edt_scan_in[106] = edt_decompressor_out[106] & bias_inputs[106];
   assign edt_scan_in[107] = edt_decompressor_out[107] & bias_inputs[107];
   assign edt_scan_in[108] = edt_decompressor_out[108] & bias_inputs[108];
   assign edt_scan_in[109] = edt_decompressor_out[109] & bias_inputs[109];
   assign edt_scan_in[110] = edt_decompressor_out[110] & bias_inputs[110];
   assign edt_scan_in[111] = edt_decompressor_out[111] & bias_inputs[111];
   assign edt_scan_in[112] = edt_decompressor_out[112] & bias_inputs[112];
   assign edt_scan_in[113] = edt_decompressor_out[113] & bias_inputs[113];
   assign edt_scan_in[114] = edt_decompressor_out[114] & bias_inputs[114];
   assign edt_scan_in[115] = edt_decompressor_out[115] & bias_inputs[115];
   assign edt_scan_in[116] = edt_decompressor_out[116] & bias_inputs[116];
   assign edt_scan_in[117] = edt_decompressor_out[117] & bias_inputs[117];
   assign edt_scan_in[118] = edt_decompressor_out[118] & bias_inputs[118];
   assign edt_scan_in[119] = edt_decompressor_out[119] & bias_inputs[119];
   assign edt_scan_in[120] = edt_decompressor_out[120] & bias_inputs[120];
   assign edt_scan_in[121] = edt_decompressor_out[121] & bias_inputs[121];
   assign edt_scan_in[122] = edt_decompressor_out[122] & bias_inputs[122];
   assign edt_scan_in[123] = edt_decompressor_out[123] & bias_inputs[123];
   assign edt_scan_in[124] = edt_decompressor_out[124] & bias_inputs[124];
   assign edt_scan_in[125] = edt_decompressor_out[125] & bias_inputs[125];
   assign edt_scan_in[126] = edt_decompressor_out[126] & bias_inputs[126];
   assign edt_scan_in[127] = edt_decompressor_out[127] & bias_inputs[127];
   assign edt_scan_in[128] = edt_decompressor_out[128] & bias_inputs[128];
   assign edt_scan_in[129] = edt_decompressor_out[129] & bias_inputs[129];
   assign edt_scan_in[130] = edt_decompressor_out[130] & bias_inputs[130];
   assign edt_scan_in[131] = edt_decompressor_out[131] & bias_inputs[131];
   assign edt_scan_in[132] = edt_decompressor_out[132] & bias_inputs[132];
   assign edt_scan_in[133] = edt_decompressor_out[133] & bias_inputs[133];
   assign edt_scan_in[134] = edt_decompressor_out[134] & bias_inputs[134];
   assign edt_scan_in[135] = edt_decompressor_out[135] & bias_inputs[135];
   assign edt_scan_in[136] = edt_decompressor_out[136] & bias_inputs[136];
   assign edt_scan_in[137] = edt_decompressor_out[137] & bias_inputs[137];
   assign edt_scan_in[138] = edt_decompressor_out[138] & bias_inputs[138];
   assign edt_scan_in[139] = edt_decompressor_out[139] & bias_inputs[139];
   assign edt_scan_in[140] = edt_decompressor_out[140] & bias_inputs[140];
   assign edt_scan_in[141] = edt_decompressor_out[141] & bias_inputs[141];
   assign edt_scan_in[142] = edt_decompressor_out[142] & bias_inputs[142];
   assign edt_scan_in[143] = edt_decompressor_out[143] & bias_inputs[143];
   assign edt_scan_in[144] = edt_decompressor_out[144] & bias_inputs[144];
   assign edt_scan_in[145] = edt_decompressor_out[145] & bias_inputs[145];
   assign edt_scan_in[146] = edt_decompressor_out[146] & bias_inputs[146];
   assign edt_scan_in[147] = edt_decompressor_out[147] & bias_inputs[147];
   assign edt_scan_in[148] = edt_decompressor_out[148] & bias_inputs[148];
   assign edt_scan_in[149] = edt_decompressor_out[149] & bias_inputs[149];
   assign edt_scan_in[150] = edt_decompressor_out[150] & bias_inputs[150];
   assign edt_scan_in[151] = edt_decompressor_out[151] & bias_inputs[151];
   assign edt_scan_in[152] = edt_decompressor_out[152] & bias_inputs[152];
   assign edt_scan_in[153] = edt_decompressor_out[153] & bias_inputs[153];
   assign edt_scan_in[154] = edt_decompressor_out[154] & bias_inputs[154];
   assign edt_scan_in[155] = edt_decompressor_out[155] & bias_inputs[155];
   assign edt_scan_in[156] = edt_decompressor_out[156] & bias_inputs[156];
   assign edt_scan_in[157] = edt_decompressor_out[157] & bias_inputs[157];
   assign edt_scan_in[158] = edt_decompressor_out[158] & bias_inputs[158];
   assign edt_scan_in[159] = edt_decompressor_out[159] & bias_inputs[159];
   assign edt_scan_in[160] = edt_decompressor_out[160] & bias_inputs[160];
   assign edt_scan_in[161] = edt_decompressor_out[161] & bias_inputs[161];
   assign edt_scan_in[162] = edt_decompressor_out[162] & bias_inputs[162];
   assign edt_scan_in[163] = edt_decompressor_out[163] & bias_inputs[163];
   assign edt_scan_in[164] = edt_decompressor_out[164] & bias_inputs[164];
   assign edt_scan_in[165] = edt_decompressor_out[165] & bias_inputs[165];
   assign edt_scan_in[166] = edt_decompressor_out[166] & bias_inputs[166];
   assign edt_scan_in[167] = edt_decompressor_out[167] & bias_inputs[167];
   assign edt_scan_in[168] = edt_decompressor_out[168] & bias_inputs[168];
   assign edt_scan_in[169] = edt_decompressor_out[169] & bias_inputs[169];
   assign edt_scan_in[170] = edt_decompressor_out[170] & bias_inputs[170];
   assign edt_scan_in[171] = edt_decompressor_out[171] & bias_inputs[171];
   assign edt_scan_in[172] = edt_decompressor_out[172] & bias_inputs[172];
   assign edt_scan_in[173] = edt_decompressor_out[173] & bias_inputs[173];
   assign edt_scan_in[174] = edt_decompressor_out[174] & bias_inputs[174];
   assign edt_scan_in[175] = edt_decompressor_out[175] & bias_inputs[175];
   assign edt_scan_in[176] = edt_decompressor_out[176] & bias_inputs[176];
   assign edt_scan_in[177] = edt_decompressor_out[177] & bias_inputs[177];
   assign edt_scan_in[178] = edt_decompressor_out[178] & bias_inputs[178];
   assign edt_scan_in[179] = edt_decompressor_out[179] & bias_inputs[179];
   assign edt_scan_in[180] = edt_decompressor_out[180] & bias_inputs[180];
   assign edt_scan_in[181] = edt_decompressor_out[181] & bias_inputs[181];
   assign edt_scan_in[182] = edt_decompressor_out[182] & bias_inputs[182];
   assign edt_scan_in[183] = edt_decompressor_out[183] & bias_inputs[183];
   assign edt_scan_in[184] = edt_decompressor_out[184] & bias_inputs[184];
   assign edt_scan_in[185] = edt_decompressor_out[185] & bias_inputs[185];
   assign edt_scan_in[186] = edt_decompressor_out[186] & bias_inputs[186];
   assign edt_scan_in[187] = edt_decompressor_out[187] & bias_inputs[187];
   assign edt_scan_in[188] = edt_decompressor_out[188] & bias_inputs[188];
   assign edt_scan_in[189] = edt_decompressor_out[189] & bias_inputs[189];
   assign edt_scan_in[190] = edt_decompressor_out[190] & bias_inputs[190];
   assign edt_scan_in[191] = edt_decompressor_out[191] & bias_inputs[191];
   assign edt_scan_in[192] = edt_decompressor_out[192] & bias_inputs[192];
   assign edt_scan_in[193] = edt_decompressor_out[193] & bias_inputs[193];
   assign edt_scan_in[194] = edt_decompressor_out[194] & bias_inputs[194];
   assign edt_scan_in[195] = edt_decompressor_out[195] & bias_inputs[195];
   assign edt_scan_in[196] = edt_decompressor_out[196] & bias_inputs[196];
   assign edt_scan_in[197] = edt_decompressor_out[197] & bias_inputs[197];
   assign edt_scan_in[198] = edt_decompressor_out[198] & bias_inputs[198];
   assign edt_scan_in[199] = edt_decompressor_out[199] & bias_inputs[199];
   assign edt_scan_in[200] = edt_decompressor_out[200] & bias_inputs[200];
   assign edt_scan_in[201] = edt_decompressor_out[201] & bias_inputs[201];
   assign edt_scan_in[202] = edt_decompressor_out[202] & bias_inputs[202];
   assign edt_scan_in[203] = edt_decompressor_out[203] & bias_inputs[203];
   assign edt_scan_in[204] = edt_decompressor_out[204] & bias_inputs[204];
   assign edt_scan_in[205] = edt_decompressor_out[205] & bias_inputs[205];
   assign edt_scan_in[206] = edt_decompressor_out[206] & bias_inputs[206];
   assign edt_scan_in[207] = edt_decompressor_out[207] & bias_inputs[207];
   assign edt_scan_in[208] = edt_decompressor_out[208] & bias_inputs[208];
   assign edt_scan_in[209] = edt_decompressor_out[209] & bias_inputs[209];
   assign edt_scan_in[210] = edt_decompressor_out[210] & bias_inputs[210];
   assign edt_scan_in[211] = edt_decompressor_out[211] & bias_inputs[211];
   assign edt_scan_in[212] = edt_decompressor_out[212] & bias_inputs[212];
   assign edt_scan_in[213] = edt_decompressor_out[213] & bias_inputs[213];
   assign edt_scan_in[214] = edt_decompressor_out[214] & bias_inputs[214];
   assign edt_scan_in[215] = edt_decompressor_out[215] & bias_inputs[215];
   assign edt_scan_in[216] = edt_decompressor_out[216] & bias_inputs[216];
   assign edt_scan_in[217] = edt_decompressor_out[217] & bias_inputs[217];
   assign edt_scan_in[218] = edt_decompressor_out[218] & bias_inputs[218];
   assign edt_scan_in[219] = edt_decompressor_out[219] & bias_inputs[219];
   assign edt_scan_in[220] = edt_decompressor_out[220] & bias_inputs[220];
   assign edt_scan_in[221] = edt_decompressor_out[221] & bias_inputs[221];
   assign edt_scan_in[222] = edt_decompressor_out[222] & bias_inputs[222];
   assign edt_scan_in[223] = edt_decompressor_out[223] & bias_inputs[223];
   assign edt_scan_in[224] = edt_decompressor_out[224] & bias_inputs[224];
   assign edt_scan_in[225] = edt_decompressor_out[225] & bias_inputs[225];
   assign edt_scan_in[226] = edt_decompressor_out[226] & bias_inputs[226];
   assign edt_scan_in[227] = edt_decompressor_out[227] & bias_inputs[227];
   assign edt_scan_in[228] = edt_decompressor_out[228] & bias_inputs[228];
   assign edt_scan_in[229] = edt_decompressor_out[229] & bias_inputs[229];
   assign edt_scan_in[230] = edt_decompressor_out[230] & bias_inputs[230];
   assign edt_scan_in[231] = edt_decompressor_out[231] & bias_inputs[231];
   assign edt_scan_in[232] = edt_decompressor_out[232] & bias_inputs[232];
   assign edt_scan_in[233] = edt_decompressor_out[233] & bias_inputs[233];
   assign edt_scan_in[234] = edt_decompressor_out[234] & bias_inputs[234];
   assign edt_scan_in[235] = edt_decompressor_out[235] & bias_inputs[235];
   assign edt_scan_in[236] = edt_decompressor_out[236] & bias_inputs[236];
   assign edt_scan_in[237] = edt_decompressor_out[237] & bias_inputs[237];
   assign edt_scan_in[238] = edt_decompressor_out[238] & bias_inputs[238];
   assign edt_scan_in[239] = edt_decompressor_out[239] & bias_inputs[239];
   assign edt_scan_in[240] = edt_decompressor_out[240] & bias_inputs[240];
   assign edt_scan_in[241] = edt_decompressor_out[241] & bias_inputs[241];
   assign edt_scan_in[242] = edt_decompressor_out[242] & bias_inputs[242];
   assign edt_scan_in[243] = edt_decompressor_out[243] & bias_inputs[243];
   assign edt_scan_in[244] = edt_decompressor_out[244] & bias_inputs[244];
   assign edt_scan_in[245] = edt_decompressor_out[245] & bias_inputs[245];
   assign edt_scan_in[246] = edt_decompressor_out[246] & bias_inputs[246];
   assign edt_scan_in[247] = edt_decompressor_out[247] & bias_inputs[247];
   assign edt_scan_in[248] = edt_decompressor_out[248] & bias_inputs[248];
   assign edt_scan_in[249] = edt_decompressor_out[249] & bias_inputs[249];
   assign edt_scan_in[250] = edt_decompressor_out[250] & bias_inputs[250];
   assign edt_scan_in[251] = edt_decompressor_out[251] & bias_inputs[251];
   assign edt_scan_in[252] = edt_decompressor_out[252] & bias_inputs[252];
   assign edt_scan_in[253] = edt_decompressor_out[253] & bias_inputs[253];
   assign edt_scan_in[254] = edt_decompressor_out[254] & bias_inputs[254];
   assign edt_scan_in[255] = edt_decompressor_out[255] & bias_inputs[255];
   assign edt_scan_in[256] = edt_decompressor_out[256] & bias_inputs[256];
   assign edt_scan_in[257] = edt_decompressor_out[257] & bias_inputs[257];
   assign edt_scan_in[258] = edt_decompressor_out[258] & bias_inputs[258];
   assign edt_scan_in[259] = edt_decompressor_out[259] & bias_inputs[259];
   assign edt_scan_in[260] = edt_decompressor_out[260] & bias_inputs[260];
   assign edt_scan_in[261] = edt_decompressor_out[261] & bias_inputs[261];
   assign edt_scan_in[262] = edt_decompressor_out[262] & bias_inputs[262];
   assign edt_scan_in[263] = edt_decompressor_out[263] & bias_inputs[263];
   assign edt_scan_in[264] = edt_decompressor_out[264] & bias_inputs[264];
   assign edt_scan_in[265] = edt_decompressor_out[265] & bias_inputs[265];
   assign edt_scan_in[266] = edt_decompressor_out[266] & bias_inputs[266];
   assign edt_scan_in[267] = edt_decompressor_out[267] & bias_inputs[267];
   assign edt_scan_in[268] = edt_decompressor_out[268] & bias_inputs[268];
   assign edt_scan_in[269] = edt_decompressor_out[269] & bias_inputs[269];
   assign edt_scan_in[270] = edt_decompressor_out[270] & bias_inputs[270];
   assign edt_scan_in[271] = edt_decompressor_out[271] & bias_inputs[271];
   assign edt_scan_in[272] = edt_decompressor_out[272] & bias_inputs[272];
   assign edt_scan_in[273] = edt_decompressor_out[273] & bias_inputs[273];
   assign edt_scan_in[274] = edt_decompressor_out[274] & bias_inputs[274];
   assign edt_scan_in[275] = edt_decompressor_out[275] & bias_inputs[275];
   assign edt_scan_in[276] = edt_decompressor_out[276] & bias_inputs[276];
   assign edt_scan_in[277] = edt_decompressor_out[277] & bias_inputs[277];
   assign edt_scan_in[278] = edt_decompressor_out[278] & bias_inputs[278];
   assign edt_scan_in[279] = edt_decompressor_out[279] & bias_inputs[279];
   assign edt_scan_in[280] = edt_decompressor_out[280] & bias_inputs[280];
   assign edt_scan_in[281] = edt_decompressor_out[281] & bias_inputs[281];
   assign edt_scan_in[282] = edt_decompressor_out[282] & bias_inputs[282];
   assign edt_scan_in[283] = edt_decompressor_out[283] & bias_inputs[283];
   assign edt_scan_in[284] = edt_decompressor_out[284] & bias_inputs[284];
   assign edt_scan_in[285] = edt_decompressor_out[285] & bias_inputs[285];
   assign edt_scan_in[286] = edt_decompressor_out[286] & bias_inputs[286];
   assign edt_scan_in[287] = edt_decompressor_out[287] & bias_inputs[287];
   assign edt_scan_in[288] = edt_decompressor_out[288] & bias_inputs[288];
   assign edt_scan_in[289] = edt_decompressor_out[289] & bias_inputs[289];
   assign edt_scan_in[290] = edt_decompressor_out[290] & bias_inputs[290];
   assign edt_scan_in[291] = edt_decompressor_out[291] & bias_inputs[291];
   assign edt_scan_in[292] = edt_decompressor_out[292] & bias_inputs[292];
   assign edt_scan_in[293] = edt_decompressor_out[293] & bias_inputs[293];
   assign edt_scan_in[294] = edt_decompressor_out[294] & bias_inputs[294];
   assign edt_scan_in[295] = edt_decompressor_out[295] & bias_inputs[295];
   assign edt_scan_in[296] = edt_decompressor_out[296] & bias_inputs[296];
   assign edt_scan_in[297] = edt_decompressor_out[297] & bias_inputs[297];
   assign edt_scan_in[298] = edt_decompressor_out[298] & bias_inputs[298];
   assign edt_scan_in[299] = edt_decompressor_out[299] & bias_inputs[299];
   assign edt_scan_in[300] = edt_decompressor_out[300] & bias_inputs[300];
   assign edt_scan_in[301] = edt_decompressor_out[301] & bias_inputs[301];
   assign edt_scan_in[302] = edt_decompressor_out[302] & bias_inputs[302];
   assign edt_scan_in[303] = edt_decompressor_out[303] & bias_inputs[303];
   assign edt_scan_in[304] = edt_decompressor_out[304] & bias_inputs[304];
   assign edt_scan_in[305] = edt_decompressor_out[305] & bias_inputs[305];
   assign edt_scan_in[306] = edt_decompressor_out[306] & bias_inputs[306];
   assign edt_scan_in[307] = edt_decompressor_out[307] & bias_inputs[307];
   assign edt_scan_in[308] = edt_decompressor_out[308] & bias_inputs[308];
   assign edt_scan_in[309] = edt_decompressor_out[309] & bias_inputs[309];
   assign edt_scan_in[310] = edt_decompressor_out[310] & bias_inputs[310];
   assign edt_scan_in[311] = edt_decompressor_out[311] & bias_inputs[311];
   assign edt_scan_in[312] = edt_decompressor_out[312] & bias_inputs[312];
   assign edt_scan_in[313] = edt_decompressor_out[313] & bias_inputs[313];
   assign edt_scan_in[314] = edt_decompressor_out[314] & bias_inputs[314];
   assign edt_scan_in[315] = edt_decompressor_out[315] & bias_inputs[315];
   assign edt_scan_in[316] = edt_decompressor_out[316] & bias_inputs[316];
   assign edt_scan_in[317] = edt_decompressor_out[317] & bias_inputs[317];
   assign edt_scan_in[318] = edt_decompressor_out[318] & bias_inputs[318];
   assign edt_scan_in[319] = edt_decompressor_out[319] & bias_inputs[319];
   assign edt_scan_in[320] = edt_decompressor_out[320] & bias_inputs[320];
   assign edt_scan_in[321] = edt_decompressor_out[321] & bias_inputs[321];
   assign edt_scan_in[322] = edt_decompressor_out[322] & bias_inputs[322];
   assign edt_scan_in[323] = edt_decompressor_out[323] & bias_inputs[323];
   assign edt_scan_in[324] = edt_decompressor_out[324] & bias_inputs[324];
   assign edt_scan_in[325] = edt_decompressor_out[325] & bias_inputs[325];
   assign edt_scan_in[326] = edt_decompressor_out[326] & bias_inputs[326];
   assign edt_scan_in[327] = edt_decompressor_out[327] & bias_inputs[327];
   assign edt_scan_in[328] = edt_decompressor_out[328] & bias_inputs[328];
   assign edt_scan_in[329] = edt_decompressor_out[329] & bias_inputs[329];
   assign edt_scan_in[330] = edt_decompressor_out[330] & bias_inputs[330];
   assign edt_scan_in[331] = edt_decompressor_out[331] & bias_inputs[331];
   assign edt_scan_in[332] = edt_decompressor_out[332] & bias_inputs[332];
   assign edt_scan_in[333] = edt_decompressor_out[333] & bias_inputs[333];
   assign edt_scan_in[334] = edt_decompressor_out[334] & bias_inputs[334];
   assign edt_scan_in[335] = edt_decompressor_out[335] & bias_inputs[335];
   assign edt_scan_in[336] = edt_decompressor_out[336] & bias_inputs[336];
   assign edt_scan_in[337] = edt_decompressor_out[337] & bias_inputs[337];
   assign edt_scan_in[338] = edt_decompressor_out[338] & bias_inputs[338];
   assign edt_scan_in[339] = edt_decompressor_out[339] & bias_inputs[339];
   assign edt_scan_in[340] = edt_decompressor_out[340] & bias_inputs[340];
   assign edt_scan_in[341] = edt_decompressor_out[341] & bias_inputs[341];
   assign edt_scan_in[342] = edt_decompressor_out[342] & bias_inputs[342];
   assign edt_scan_in[343] = edt_decompressor_out[343] & bias_inputs[343];
   assign edt_scan_in[344] = edt_decompressor_out[344] & bias_inputs[344];
   assign edt_scan_in[345] = edt_decompressor_out[345] & bias_inputs[345];
   assign edt_scan_in[346] = edt_decompressor_out[346] & bias_inputs[346];
   assign edt_scan_in[347] = edt_decompressor_out[347] & bias_inputs[347];
   assign edt_scan_in[348] = edt_decompressor_out[348] & bias_inputs[348];
   assign edt_scan_in[349] = edt_decompressor_out[349] & bias_inputs[349];
   assign edt_scan_in[350] = edt_decompressor_out[350] & bias_inputs[350];
   assign edt_scan_in[351] = edt_decompressor_out[351] & bias_inputs[351];
   assign edt_scan_in[352] = edt_decompressor_out[352] & bias_inputs[352];
   assign edt_scan_in[353] = edt_decompressor_out[353] & bias_inputs[353];
   assign edt_scan_in[354] = edt_decompressor_out[354] & bias_inputs[354];
   assign edt_scan_in[355] = edt_decompressor_out[355] & bias_inputs[355];
   assign edt_scan_in[356] = edt_decompressor_out[356] & bias_inputs[356];
   assign edt_scan_in[357] = edt_decompressor_out[357] & bias_inputs[357];
   assign edt_scan_in[358] = edt_decompressor_out[358] & bias_inputs[358];
   assign edt_scan_in[359] = edt_decompressor_out[359] & bias_inputs[359];
   assign edt_scan_in[360] = edt_decompressor_out[360] & bias_inputs[360];
   assign edt_scan_in[361] = edt_decompressor_out[361] & bias_inputs[361];
   assign edt_scan_in[362] = edt_decompressor_out[362] & bias_inputs[362];
   assign edt_scan_in[363] = edt_decompressor_out[363] & bias_inputs[363];
   assign edt_scan_in[364] = edt_decompressor_out[364] & bias_inputs[364];
   assign edt_scan_in[365] = edt_decompressor_out[365] & bias_inputs[365];
   assign edt_scan_in[366] = edt_decompressor_out[366] & bias_inputs[366];
   assign edt_scan_in[367] = edt_decompressor_out[367] & bias_inputs[367];
   assign edt_scan_in[368] = edt_decompressor_out[368] & bias_inputs[368];
   assign edt_scan_in[369] = edt_decompressor_out[369] & bias_inputs[369];
   assign edt_scan_in[370] = edt_decompressor_out[370] & bias_inputs[370];
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_onehot_decoder_8_to_185 (
   input  wire [  7:0] encoded_masks,
   output reg  [184:0] decoded_masks
);
   always @(encoded_masks)
   begin
      case (encoded_masks)
         8'b00000000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b00000001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
         8'b00000010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
         8'b00000011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
         8'b00000100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
         8'b00000101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
         8'b00000110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
         8'b00000111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
         8'b00001000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
         8'b00001001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
         8'b00001010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
         8'b00001011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
         8'b00001100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
         8'b00001101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
         8'b00001110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
         8'b00001111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
         8'b00010000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
         8'b00010001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
         8'b00010010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
         8'b00010011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
         8'b00010100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
         8'b00010101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
         8'b00010110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
         8'b00010111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
         8'b00011000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
         8'b00011001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
         8'b00011010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
         8'b00011011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
         8'b00011100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
         8'b00011101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
         8'b00011110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
         8'b00011111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
         8'b00100000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
         8'b00100001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
         8'b00100010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
         8'b00100011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
         8'b00100100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
         8'b00100101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
         8'b00100110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
         8'b00100111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
         8'b00101000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
         8'b00101001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
         8'b00101010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
         8'b00101011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
         8'b00101100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
         8'b00101101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
         8'b00101110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
         8'b00101111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
         8'b00110000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
         8'b00110001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
         8'b00110010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
         8'b00110011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
         8'b00110100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
         8'b00110101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
         8'b00110110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
         8'b00110111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
         8'b00111000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
         8'b00111001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
         8'b00111010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
         8'b00111011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
         8'b00111100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
         8'b00111101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
         8'b00111110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
         8'b00111111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
         8'b01000000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
         8'b01000001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
         8'b01000010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
         8'b01000011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000000: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000001: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000010: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000011: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000100: decoded_masks = 185'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000101: decoded_masks = 185'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000110: decoded_masks = 185'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000111: decoded_masks = 185'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001000: decoded_masks = 185'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001001: decoded_masks = 185'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001010: decoded_masks = 185'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001011: decoded_masks = 185'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001100: decoded_masks = 185'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001101: decoded_masks = 185'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001110: decoded_masks = 185'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001111: decoded_masks = 185'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010000: decoded_masks = 185'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010001: decoded_masks = 185'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010010: decoded_masks = 185'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010011: decoded_masks = 185'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010100: decoded_masks = 185'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010101: decoded_masks = 185'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010110: decoded_masks = 185'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010111: decoded_masks = 185'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011000: decoded_masks = 185'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011001: decoded_masks = 185'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011010: decoded_masks = 185'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011011: decoded_masks = 185'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011100: decoded_masks = 185'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011101: decoded_masks = 185'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011110: decoded_masks = 185'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011111: decoded_masks = 185'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100000: decoded_masks = 185'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100001: decoded_masks = 185'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100010: decoded_masks = 185'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100011: decoded_masks = 185'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100100: decoded_masks = 185'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100101: decoded_masks = 185'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100110: decoded_masks = 185'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100111: decoded_masks = 185'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101000: decoded_masks = 185'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101001: decoded_masks = 185'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101010: decoded_masks = 185'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101011: decoded_masks = 185'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101100: decoded_masks = 185'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101101: decoded_masks = 185'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101110: decoded_masks = 185'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101111: decoded_masks = 185'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110000: decoded_masks = 185'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110001: decoded_masks = 185'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110010: decoded_masks = 185'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110011: decoded_masks = 185'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110100: decoded_masks = 185'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110101: decoded_masks = 185'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110110: decoded_masks = 185'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110111: decoded_masks = 185'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10111000: decoded_masks = 185'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10111001: decoded_masks = 185'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         default:     decoded_masks = 185'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
      endcase
   end
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_onehot_decoder_8_to_186 (
   input  wire [  7:0] encoded_masks,
   output reg  [185:0] decoded_masks
);
   always @(encoded_masks)
   begin
      case (encoded_masks)
         8'b00000000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b00000001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
         8'b00000010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
         8'b00000011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
         8'b00000100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
         8'b00000101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
         8'b00000110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
         8'b00000111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
         8'b00001000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
         8'b00001001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
         8'b00001010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
         8'b00001011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
         8'b00001100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
         8'b00001101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
         8'b00001110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
         8'b00001111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
         8'b00010000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
         8'b00010001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
         8'b00010010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
         8'b00010011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
         8'b00010100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
         8'b00010101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
         8'b00010110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
         8'b00010111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
         8'b00011000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
         8'b00011001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
         8'b00011010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
         8'b00011011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
         8'b00011100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
         8'b00011101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
         8'b00011110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
         8'b00011111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
         8'b00100000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
         8'b00100001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
         8'b00100010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
         8'b00100011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
         8'b00100100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
         8'b00100101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
         8'b00100110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
         8'b00100111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
         8'b00101000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
         8'b00101001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
         8'b00101010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
         8'b00101011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
         8'b00101100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
         8'b00101101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
         8'b00101110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
         8'b00101111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
         8'b00110000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
         8'b00110001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
         8'b00110010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
         8'b00110011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
         8'b00110100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
         8'b00110101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
         8'b00110110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
         8'b00110111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
         8'b00111000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
         8'b00111001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
         8'b00111010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
         8'b00111011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
         8'b00111100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
         8'b00111101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
         8'b00111110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
         8'b00111111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
         8'b01000000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
         8'b01000001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
         8'b01000010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
         8'b01000011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01000111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01001111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01010111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01011111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01100111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01101111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01110111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b01111111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000000: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000001: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000010: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000011: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000100: decoded_masks = 186'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000101: decoded_masks = 186'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000110: decoded_masks = 186'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10000111: decoded_masks = 186'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001000: decoded_masks = 186'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001001: decoded_masks = 186'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001010: decoded_masks = 186'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001011: decoded_masks = 186'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001100: decoded_masks = 186'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001101: decoded_masks = 186'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001110: decoded_masks = 186'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10001111: decoded_masks = 186'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010000: decoded_masks = 186'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010001: decoded_masks = 186'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010010: decoded_masks = 186'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010011: decoded_masks = 186'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010100: decoded_masks = 186'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010101: decoded_masks = 186'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010110: decoded_masks = 186'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10010111: decoded_masks = 186'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011000: decoded_masks = 186'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011001: decoded_masks = 186'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011010: decoded_masks = 186'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011011: decoded_masks = 186'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011100: decoded_masks = 186'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011101: decoded_masks = 186'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011110: decoded_masks = 186'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10011111: decoded_masks = 186'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100000: decoded_masks = 186'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100001: decoded_masks = 186'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100010: decoded_masks = 186'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100011: decoded_masks = 186'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100100: decoded_masks = 186'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100101: decoded_masks = 186'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100110: decoded_masks = 186'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10100111: decoded_masks = 186'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101000: decoded_masks = 186'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101001: decoded_masks = 186'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101010: decoded_masks = 186'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101011: decoded_masks = 186'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101100: decoded_masks = 186'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101101: decoded_masks = 186'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101110: decoded_masks = 186'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10101111: decoded_masks = 186'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110000: decoded_masks = 186'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110001: decoded_masks = 186'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110010: decoded_masks = 186'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110011: decoded_masks = 186'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110100: decoded_masks = 186'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110101: decoded_masks = 186'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110110: decoded_masks = 186'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10110111: decoded_masks = 186'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10111000: decoded_masks = 186'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10111001: decoded_masks = 186'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         8'b10111010: decoded_masks = 186'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
         default:     decoded_masks = 186'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
      endcase
   end
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_xor_decoder (
   input  wire [ 29:0] encoded_masks,
   output wire [185:0] decoded_masks_0,
   output wire [184:0] decoded_masks_1
);
   assign decoded_masks_0[  0] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 2];
   assign decoded_masks_0[  1] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 3];
   assign decoded_masks_0[  2] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 4];
   assign decoded_masks_0[  3] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 5];
   assign decoded_masks_0[  4] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 6];
   assign decoded_masks_0[  5] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 7];
   assign decoded_masks_0[  6] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 8];
   assign decoded_masks_0[  7] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[ 9];
   assign decoded_masks_0[  8] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[10];
   assign decoded_masks_0[  9] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[11];
   assign decoded_masks_0[ 10] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[12];
   assign decoded_masks_0[ 11] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[13];
   assign decoded_masks_0[ 12] = encoded_masks[ 0] ^ encoded_masks[ 1] ^ encoded_masks[14];
   assign decoded_masks_0[ 13] = encoded_masks[ 0] ^ encoded_masks[ 2] ^ encoded_masks[ 3];
   assign decoded_masks_0[ 14] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[ 3];
   assign decoded_masks_0[ 15] = encoded_masks[ 8] ^ encoded_masks[11] ^ encoded_masks[13];
   assign decoded_masks_0[ 16] = encoded_masks[ 0] ^ encoded_masks[ 9] ^ encoded_masks[12];
   assign decoded_masks_0[ 17] = encoded_masks[ 4] ^ encoded_masks[ 6] ^ encoded_masks[ 7];
   assign decoded_masks_0[ 18] = encoded_masks[ 5] ^ encoded_masks[10] ^ encoded_masks[14];
   assign decoded_masks_0[ 19] = encoded_masks[ 1] ^ encoded_masks[ 5] ^ encoded_masks[13];
   assign decoded_masks_0[ 20] = encoded_masks[ 4] ^ encoded_masks[ 8] ^ encoded_masks[12];
   assign decoded_masks_0[ 21] = encoded_masks[ 3] ^ encoded_masks[ 7] ^ encoded_masks[10];
   assign decoded_masks_0[ 22] = encoded_masks[ 6] ^ encoded_masks[ 9] ^ encoded_masks[14];
   assign decoded_masks_0[ 23] = encoded_masks[ 2] ^ encoded_masks[ 6] ^ encoded_masks[11];
   assign decoded_masks_0[ 24] = encoded_masks[10] ^ encoded_masks[11] ^ encoded_masks[12];
   assign decoded_masks_0[ 25] = encoded_masks[ 5] ^ encoded_masks[ 7] ^ encoded_masks[ 8];
   assign decoded_masks_0[ 26] = encoded_masks[ 0] ^ encoded_masks[ 4] ^ encoded_masks[14];
   assign decoded_masks_0[ 27] = encoded_masks[ 3] ^ encoded_masks[ 9] ^ encoded_masks[13];
   assign decoded_masks_0[ 28] = encoded_masks[ 2] ^ encoded_masks[ 8] ^ encoded_masks[10];
   assign decoded_masks_0[ 29] = encoded_masks[ 4] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[ 30] = encoded_masks[ 7] ^ encoded_masks[12] ^ encoded_masks[13];
   assign decoded_masks_0[ 31] = encoded_masks[ 3] ^ encoded_masks[ 5] ^ encoded_masks[ 6];
   assign decoded_masks_0[ 32] = encoded_masks[ 2] ^ encoded_masks[12] ^ encoded_masks[14];
   assign decoded_masks_0[ 33] = encoded_masks[ 1] ^ encoded_masks[ 8] ^ encoded_masks[11];
   assign decoded_masks_0[ 34] = encoded_masks[ 0] ^ encoded_masks[ 6] ^ encoded_masks[ 7];
   assign decoded_masks_0[ 35] = encoded_masks[ 9] ^ encoded_masks[10] ^ encoded_masks[13];
   assign decoded_masks_0[ 36] = encoded_masks[ 2] ^ encoded_masks[ 4] ^ encoded_masks[ 5];
   assign decoded_masks_0[ 37] = encoded_masks[ 3] ^ encoded_masks[11] ^ encoded_masks[14];
   assign decoded_masks_0[ 38] = encoded_masks[ 7] ^ encoded_masks[ 9] ^ encoded_masks[14];
   assign decoded_masks_0[ 39] = encoded_masks[ 4] ^ encoded_masks[ 6] ^ encoded_masks[13];
   assign decoded_masks_0[ 40] = encoded_masks[ 3] ^ encoded_masks[ 8] ^ encoded_masks[12];
   assign decoded_masks_0[ 41] = encoded_masks[ 5] ^ encoded_masks[ 8] ^ encoded_masks[ 9];
   assign decoded_masks_0[ 42] = encoded_masks[ 1] ^ encoded_masks[10] ^ encoded_masks[14];
   assign decoded_masks_0[ 43] = encoded_masks[ 6] ^ encoded_masks[10] ^ encoded_masks[12];
   assign decoded_masks_0[ 44] = encoded_masks[ 2] ^ encoded_masks[ 7] ^ encoded_masks[13];
   assign decoded_masks_0[ 45] = encoded_masks[ 4] ^ encoded_masks[ 5] ^ encoded_masks[11];
   assign decoded_masks_0[ 46] = encoded_masks[ 1] ^ encoded_masks[ 5] ^ encoded_masks[ 9];
   assign decoded_masks_0[ 47] = encoded_masks[ 8] ^ encoded_masks[13] ^ encoded_masks[14];
   assign decoded_masks_0[ 48] = encoded_masks[ 3] ^ encoded_masks[ 7] ^ encoded_masks[12];
   assign decoded_masks_0[ 49] = encoded_masks[ 0] ^ encoded_masks[ 4] ^ encoded_masks[10];
   assign decoded_masks_0[ 50] = encoded_masks[ 3] ^ encoded_masks[ 6] ^ encoded_masks[11];
   assign decoded_masks_0[ 51] = encoded_masks[ 2] ^ encoded_masks[ 4] ^ encoded_masks[12];
   assign decoded_masks_0[ 52] = encoded_masks[ 6] ^ encoded_masks[ 8] ^ encoded_masks[14];
   assign decoded_masks_0[ 53] = encoded_masks[ 2] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[ 54] = encoded_masks[ 7] ^ encoded_masks[11] ^ encoded_masks[14];
   assign decoded_masks_0[ 55] = encoded_masks[ 2] ^ encoded_masks[10] ^ encoded_masks[13];
   assign decoded_masks_0[ 56] = encoded_masks[ 1] ^ encoded_masks[ 5] ^ encoded_masks[12];
   assign decoded_masks_0[ 57] = encoded_masks[ 3] ^ encoded_masks[ 4] ^ encoded_masks[ 5];
   assign decoded_masks_0[ 58] = encoded_masks[ 8] ^ encoded_masks[ 9] ^ encoded_masks[10];
   assign decoded_masks_0[ 59] = encoded_masks[ 6] ^ encoded_masks[ 7] ^ encoded_masks[13];
   assign decoded_masks_0[ 60] = encoded_masks[ 5] ^ encoded_masks[ 7] ^ encoded_masks[10];
   assign decoded_masks_0[ 61] = encoded_masks[ 2] ^ encoded_masks[ 6] ^ encoded_masks[ 8];
   assign decoded_masks_0[ 62] = encoded_masks[ 0] ^ encoded_masks[ 9] ^ encoded_masks[13];
   assign decoded_masks_0[ 63] = encoded_masks[11] ^ encoded_masks[12] ^ encoded_masks[14];
   assign decoded_masks_0[ 64] = encoded_masks[ 3] ^ encoded_masks[ 5] ^ encoded_masks[ 8];
   assign decoded_masks_0[ 65] = encoded_masks[ 3] ^ encoded_masks[ 4] ^ encoded_masks[ 7];
   assign decoded_masks_0[ 66] = encoded_masks[ 0] ^ encoded_masks[ 9] ^ encoded_masks[14];
   assign decoded_masks_0[ 67] = encoded_masks[ 4] ^ encoded_masks[ 6] ^ encoded_masks[10];
   assign decoded_masks_0[ 68] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[13];
   assign decoded_masks_0[ 69] = encoded_masks[ 5] ^ encoded_masks[ 6] ^ encoded_masks[12];
   assign decoded_masks_0[ 70] = encoded_masks[ 2] ^ encoded_masks[ 8] ^ encoded_masks[11];
   assign decoded_masks_0[ 71] = encoded_masks[ 4] ^ encoded_masks[12] ^ encoded_masks[14];
   assign decoded_masks_0[ 72] = encoded_masks[ 0] ^ encoded_masks[ 3] ^ encoded_masks[ 7];
   assign decoded_masks_0[ 73] = encoded_masks[ 5] ^ encoded_masks[ 9] ^ encoded_masks[10];
   assign decoded_masks_0[ 74] = encoded_masks[ 0] ^ encoded_masks[ 6] ^ encoded_masks[11];
   assign decoded_masks_0[ 75] = encoded_masks[ 3] ^ encoded_masks[11] ^ encoded_masks[13];
   assign decoded_masks_0[ 76] = encoded_masks[ 7] ^ encoded_masks[ 9] ^ encoded_masks[12];
   assign decoded_masks_0[ 77] = encoded_masks[ 4] ^ encoded_masks[10] ^ encoded_masks[14];
   assign decoded_masks_0[ 78] = encoded_masks[ 3] ^ encoded_masks[ 8] ^ encoded_masks[ 9];
   assign decoded_masks_0[ 79] = encoded_masks[10] ^ encoded_masks[13] ^ encoded_masks[14];
   assign decoded_masks_0[ 80] = encoded_masks[ 2] ^ encoded_masks[ 5] ^ encoded_masks[ 6];
   assign decoded_masks_0[ 81] = encoded_masks[ 1] ^ encoded_masks[ 7] ^ encoded_masks[ 8];
   assign decoded_masks_0[ 82] = encoded_masks[ 5] ^ encoded_masks[11] ^ encoded_masks[12];
   assign decoded_masks_0[ 83] = encoded_masks[ 0] ^ encoded_masks[ 4] ^ encoded_masks[11];
   assign decoded_masks_0[ 84] = encoded_masks[ 2] ^ encoded_masks[ 4] ^ encoded_masks[ 7];
   assign decoded_masks_0[ 85] = encoded_masks[ 9] ^ encoded_masks[13] ^ encoded_masks[14];
   assign decoded_masks_0[ 86] = encoded_masks[ 1] ^ encoded_masks[ 6] ^ encoded_masks[10];
   assign decoded_masks_0[ 87] = encoded_masks[ 2] ^ encoded_masks[ 3] ^ encoded_masks[12];
   assign decoded_masks_0[ 88] = encoded_masks[ 4] ^ encoded_masks[ 9] ^ encoded_masks[13];
   assign decoded_masks_0[ 89] = encoded_masks[ 3] ^ encoded_masks[10] ^ encoded_masks[12];
   assign decoded_masks_0[ 90] = encoded_masks[ 5] ^ encoded_masks[ 8] ^ encoded_masks[13];
   assign decoded_masks_0[ 91] = encoded_masks[ 7] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[ 92] = encoded_masks[ 4] ^ encoded_masks[ 6] ^ encoded_masks[ 8];
   assign decoded_masks_0[ 93] = encoded_masks[ 0] ^ encoded_masks[ 2] ^ encoded_masks[14];
   assign decoded_masks_0[ 94] = encoded_masks[ 1] ^ encoded_masks[ 6] ^ encoded_masks[13];
   assign decoded_masks_0[ 95] = encoded_masks[ 8] ^ encoded_masks[10] ^ encoded_masks[14];
   assign decoded_masks_0[ 96] = encoded_masks[ 5] ^ encoded_masks[ 7] ^ encoded_masks[11];
   assign decoded_masks_0[ 97] = encoded_masks[ 2] ^ encoded_masks[ 3] ^ encoded_masks[ 9];
   assign decoded_masks_0[ 98] = encoded_masks[ 0] ^ encoded_masks[ 5] ^ encoded_masks[12];
   assign decoded_masks_0[ 99] = encoded_masks[ 3] ^ encoded_masks[ 8] ^ encoded_masks[10];
   assign decoded_masks_0[100] = encoded_masks[12] ^ encoded_masks[13] ^ encoded_masks[14];
   assign decoded_masks_0[101] = encoded_masks[ 4] ^ encoded_masks[ 5] ^ encoded_masks[ 7];
   assign decoded_masks_0[102] = encoded_masks[ 2] ^ encoded_masks[11] ^ encoded_masks[12];
   assign decoded_masks_0[103] = encoded_masks[ 1] ^ encoded_masks[ 4] ^ encoded_masks[10];
   assign decoded_masks_0[104] = encoded_masks[ 2] ^ encoded_masks[ 6] ^ encoded_masks[ 9];
   assign decoded_masks_0[105] = encoded_masks[ 7] ^ encoded_masks[10] ^ encoded_masks[11];
   assign decoded_masks_0[106] = encoded_masks[ 0] ^ encoded_masks[ 6] ^ encoded_masks[13];
   assign decoded_masks_0[107] = encoded_masks[ 3] ^ encoded_masks[ 4] ^ encoded_masks[14];
   assign decoded_masks_0[108] = encoded_masks[ 8] ^ encoded_masks[12] ^ encoded_masks[13];
   assign decoded_masks_0[109] = encoded_masks[ 1] ^ encoded_masks[ 7] ^ encoded_masks[11];
   assign decoded_masks_0[110] = encoded_masks[ 5] ^ encoded_masks[12] ^ encoded_masks[14];
   assign decoded_masks_0[111] = encoded_masks[ 5] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[112] = encoded_masks[ 0] ^ encoded_masks[ 7] ^ encoded_masks[ 8];
   assign decoded_masks_0[113] = encoded_masks[ 2] ^ encoded_masks[ 6] ^ encoded_masks[14];
   assign decoded_masks_0[114] = encoded_masks[ 2] ^ encoded_masks[ 3] ^ encoded_masks[13];
   assign decoded_masks_0[115] = encoded_masks[ 3] ^ encoded_masks[ 4] ^ encoded_masks[10];
   assign decoded_masks_0[116] = encoded_masks[ 0] ^ encoded_masks[ 8] ^ encoded_masks[11];
   assign decoded_masks_0[117] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[14];
   assign decoded_masks_0[118] = encoded_masks[ 6] ^ encoded_masks[ 8] ^ encoded_masks[12];
   assign decoded_masks_0[119] = encoded_masks[ 4] ^ encoded_masks[ 5] ^ encoded_masks[13];
   assign decoded_masks_0[120] = encoded_masks[ 2] ^ encoded_masks[ 9] ^ encoded_masks[10];
   assign decoded_masks_0[121] = encoded_masks[ 3] ^ encoded_masks[ 6] ^ encoded_masks[14];
   assign decoded_masks_0[122] = encoded_masks[ 4] ^ encoded_masks[ 8] ^ encoded_masks[ 9];
   assign decoded_masks_0[123] = encoded_masks[ 0] ^ encoded_masks[ 7] ^ encoded_masks[10];
   assign decoded_masks_0[124] = encoded_masks[ 3] ^ encoded_masks[ 6] ^ encoded_masks[12];
   assign decoded_masks_0[125] = encoded_masks[ 7] ^ encoded_masks[ 8] ^ encoded_masks[13];
   assign decoded_masks_0[126] = encoded_masks[ 1] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[127] = encoded_masks[ 5] ^ encoded_masks[11] ^ encoded_masks[13];
   assign decoded_masks_0[128] = encoded_masks[ 2] ^ encoded_masks[ 7] ^ encoded_masks[14];
   assign decoded_masks_0[129] = encoded_masks[ 1] ^ encoded_masks[ 3] ^ encoded_masks[10];
   assign decoded_masks_0[130] = encoded_masks[ 1] ^ encoded_masks[ 3] ^ encoded_masks[ 4];
   assign decoded_masks_0[131] = encoded_masks[ 6] ^ encoded_masks[ 9] ^ encoded_masks[11];
   assign decoded_masks_0[132] = encoded_masks[ 2] ^ encoded_masks[ 8] ^ encoded_masks[12];
   assign decoded_masks_0[133] = encoded_masks[ 0] ^ encoded_masks[ 5] ^ encoded_masks[13];
   assign decoded_masks_0[134] = encoded_masks[ 4] ^ encoded_masks[ 9] ^ encoded_masks[14];
   assign decoded_masks_0[135] = encoded_masks[ 0] ^ encoded_masks[ 5] ^ encoded_masks[ 6];
   assign decoded_masks_0[136] = encoded_masks[ 7] ^ encoded_masks[ 8] ^ encoded_masks[10];
   assign decoded_masks_0[137] = encoded_masks[10] ^ encoded_masks[12] ^ encoded_masks[13];
   assign decoded_masks_0[138] = encoded_masks[ 4] ^ encoded_masks[ 6] ^ encoded_masks[14];
   assign decoded_masks_0[139] = encoded_masks[ 1] ^ encoded_masks[ 7] ^ encoded_masks[ 9];
   assign decoded_masks_0[140] = encoded_masks[ 5] ^ encoded_masks[13] ^ encoded_masks[14];
   assign decoded_masks_0[141] = encoded_masks[ 4] ^ encoded_masks[11] ^ encoded_masks[12];
   assign decoded_masks_0[142] = encoded_masks[ 1] ^ encoded_masks[ 3] ^ encoded_masks[12];
   assign decoded_masks_0[143] = encoded_masks[ 2] ^ encoded_masks[ 3] ^ encoded_masks[11];
   assign decoded_masks_0[144] = encoded_masks[ 2] ^ encoded_masks[ 5] ^ encoded_masks[ 7];
   assign decoded_masks_0[145] = encoded_masks[ 0] ^ encoded_masks[ 6] ^ encoded_masks[10];
   assign decoded_masks_0[146] = encoded_masks[ 5] ^ encoded_masks[ 8] ^ encoded_masks[14];
   assign decoded_masks_0[147] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[ 9];
   assign decoded_masks_0[148] = encoded_masks[ 3] ^ encoded_masks[ 6] ^ encoded_masks[13];
   assign decoded_masks_0[149] = encoded_masks[ 7] ^ encoded_masks[ 8] ^ encoded_masks[ 9];
   assign decoded_masks_0[150] = encoded_masks[ 7] ^ encoded_masks[11] ^ encoded_masks[13];
   assign decoded_masks_0[151] = encoded_masks[ 5] ^ encoded_masks[11] ^ encoded_masks[14];
   assign decoded_masks_0[152] = encoded_masks[ 4] ^ encoded_masks[10] ^ encoded_masks[12];
   assign decoded_masks_0[153] = encoded_masks[ 0] ^ encoded_masks[ 3] ^ encoded_masks[ 8];
   assign decoded_masks_0[154] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[ 4];
   assign decoded_masks_0[155] = encoded_masks[ 6] ^ encoded_masks[ 9] ^ encoded_masks[12];
   assign decoded_masks_0[156] = encoded_masks[ 3] ^ encoded_masks[ 7] ^ encoded_masks[14];
   assign decoded_masks_0[157] = encoded_masks[ 7] ^ encoded_masks[ 9] ^ encoded_masks[10];
   assign decoded_masks_0[158] = encoded_masks[ 4] ^ encoded_masks[ 5] ^ encoded_masks[ 8];
   assign decoded_masks_0[159] = encoded_masks[ 0] ^ encoded_masks[11] ^ encoded_masks[12];
   assign decoded_masks_0[160] = encoded_masks[ 1] ^ encoded_masks[ 6] ^ encoded_masks[12];
   assign decoded_masks_0[161] = encoded_masks[10] ^ encoded_masks[11] ^ encoded_masks[13];
   assign decoded_masks_0[162] = encoded_masks[ 2] ^ encoded_masks[ 3] ^ encoded_masks[ 4];
   assign decoded_masks_0[163] = encoded_masks[ 6] ^ encoded_masks[ 9] ^ encoded_masks[13];
   assign decoded_masks_0[164] = encoded_masks[ 1] ^ encoded_masks[ 2] ^ encoded_masks[ 8];
   assign decoded_masks_0[165] = encoded_masks[ 2] ^ encoded_masks[ 5] ^ encoded_masks[10];
   assign decoded_masks_0[166] = encoded_masks[ 5] ^ encoded_masks[10] ^ encoded_masks[11];
   assign decoded_masks_0[167] = encoded_masks[ 3] ^ encoded_masks[ 9] ^ encoded_masks[14];
   assign decoded_masks_0[168] = encoded_masks[ 4] ^ encoded_masks[ 8] ^ encoded_masks[11];
   assign decoded_masks_0[169] = encoded_masks[ 7] ^ encoded_masks[10] ^ encoded_masks[12];
   assign decoded_masks_0[170] = encoded_masks[ 6] ^ encoded_masks[12] ^ encoded_masks[14];
   assign decoded_masks_0[171] = encoded_masks[ 0] ^ encoded_masks[ 4] ^ encoded_masks[ 9];
   assign decoded_masks_0[172] = encoded_masks[ 2] ^ encoded_masks[ 5] ^ encoded_masks[12];
   assign decoded_masks_0[173] = encoded_masks[ 1] ^ encoded_masks[ 6] ^ encoded_masks[ 7];
   assign decoded_masks_0[174] = encoded_masks[ 1] ^ encoded_masks[ 8] ^ encoded_masks[14];
   assign decoded_masks_0[175] = encoded_masks[ 0] ^ encoded_masks[ 2] ^ encoded_masks[13];
   assign decoded_masks_0[176] = encoded_masks[ 3] ^ encoded_masks[ 5] ^ encoded_masks[ 9];
   assign decoded_masks_0[177] = encoded_masks[ 0] ^ encoded_masks[ 4] ^ encoded_masks[13];
   assign decoded_masks_0[178] = encoded_masks[ 1] ^ encoded_masks[ 7] ^ encoded_masks[12];
   assign decoded_masks_0[179] = encoded_masks[ 0] ^ encoded_masks[ 3] ^ encoded_masks[14];
   assign decoded_masks_0[180] = encoded_masks[ 6] ^ encoded_masks[ 8] ^ encoded_masks[13];
   assign decoded_masks_0[181] = encoded_masks[ 2] ^ encoded_masks[ 6] ^ encoded_masks[10];
   assign decoded_masks_0[182] = encoded_masks[ 2] ^ encoded_masks[ 4] ^ encoded_masks[11];
   assign decoded_masks_0[183] = encoded_masks[ 5] ^ encoded_masks[ 9] ^ encoded_masks[13];
   assign decoded_masks_0[184] = encoded_masks[ 8] ^ encoded_masks[10] ^ encoded_masks[11];
   assign decoded_masks_0[185] = encoded_masks[ 0] ^ encoded_masks[ 8] ^ encoded_masks[12];

   assign decoded_masks_1[  0] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[17];
   assign decoded_masks_1[  1] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[18];
   assign decoded_masks_1[  2] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[19];
   assign decoded_masks_1[  3] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[20];
   assign decoded_masks_1[  4] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[21];
   assign decoded_masks_1[  5] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[22];
   assign decoded_masks_1[  6] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[23];
   assign decoded_masks_1[  7] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[24];
   assign decoded_masks_1[  8] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[25];
   assign decoded_masks_1[  9] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[26];
   assign decoded_masks_1[ 10] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[27];
   assign decoded_masks_1[ 11] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[28];
   assign decoded_masks_1[ 12] = encoded_masks[15] ^ encoded_masks[16] ^ encoded_masks[29];
   assign decoded_masks_1[ 13] = encoded_masks[15] ^ encoded_masks[17] ^ encoded_masks[18];
   assign decoded_masks_1[ 14] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[18];
   assign decoded_masks_1[ 15] = encoded_masks[23] ^ encoded_masks[26] ^ encoded_masks[28];
   assign decoded_masks_1[ 16] = encoded_masks[15] ^ encoded_masks[24] ^ encoded_masks[27];
   assign decoded_masks_1[ 17] = encoded_masks[19] ^ encoded_masks[21] ^ encoded_masks[22];
   assign decoded_masks_1[ 18] = encoded_masks[20] ^ encoded_masks[25] ^ encoded_masks[29];
   assign decoded_masks_1[ 19] = encoded_masks[16] ^ encoded_masks[20] ^ encoded_masks[28];
   assign decoded_masks_1[ 20] = encoded_masks[19] ^ encoded_masks[23] ^ encoded_masks[27];
   assign decoded_masks_1[ 21] = encoded_masks[18] ^ encoded_masks[22] ^ encoded_masks[25];
   assign decoded_masks_1[ 22] = encoded_masks[21] ^ encoded_masks[24] ^ encoded_masks[29];
   assign decoded_masks_1[ 23] = encoded_masks[17] ^ encoded_masks[21] ^ encoded_masks[26];
   assign decoded_masks_1[ 24] = encoded_masks[25] ^ encoded_masks[26] ^ encoded_masks[27];
   assign decoded_masks_1[ 25] = encoded_masks[20] ^ encoded_masks[22] ^ encoded_masks[23];
   assign decoded_masks_1[ 26] = encoded_masks[15] ^ encoded_masks[19] ^ encoded_masks[29];
   assign decoded_masks_1[ 27] = encoded_masks[18] ^ encoded_masks[24] ^ encoded_masks[28];
   assign decoded_masks_1[ 28] = encoded_masks[17] ^ encoded_masks[23] ^ encoded_masks[25];
   assign decoded_masks_1[ 29] = encoded_masks[19] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[ 30] = encoded_masks[22] ^ encoded_masks[27] ^ encoded_masks[28];
   assign decoded_masks_1[ 31] = encoded_masks[18] ^ encoded_masks[20] ^ encoded_masks[21];
   assign decoded_masks_1[ 32] = encoded_masks[17] ^ encoded_masks[27] ^ encoded_masks[29];
   assign decoded_masks_1[ 33] = encoded_masks[16] ^ encoded_masks[23] ^ encoded_masks[26];
   assign decoded_masks_1[ 34] = encoded_masks[15] ^ encoded_masks[21] ^ encoded_masks[22];
   assign decoded_masks_1[ 35] = encoded_masks[24] ^ encoded_masks[25] ^ encoded_masks[28];
   assign decoded_masks_1[ 36] = encoded_masks[17] ^ encoded_masks[19] ^ encoded_masks[20];
   assign decoded_masks_1[ 37] = encoded_masks[18] ^ encoded_masks[26] ^ encoded_masks[29];
   assign decoded_masks_1[ 38] = encoded_masks[22] ^ encoded_masks[24] ^ encoded_masks[29];
   assign decoded_masks_1[ 39] = encoded_masks[19] ^ encoded_masks[21] ^ encoded_masks[28];
   assign decoded_masks_1[ 40] = encoded_masks[18] ^ encoded_masks[23] ^ encoded_masks[27];
   assign decoded_masks_1[ 41] = encoded_masks[20] ^ encoded_masks[23] ^ encoded_masks[24];
   assign decoded_masks_1[ 42] = encoded_masks[16] ^ encoded_masks[25] ^ encoded_masks[29];
   assign decoded_masks_1[ 43] = encoded_masks[21] ^ encoded_masks[25] ^ encoded_masks[27];
   assign decoded_masks_1[ 44] = encoded_masks[17] ^ encoded_masks[22] ^ encoded_masks[28];
   assign decoded_masks_1[ 45] = encoded_masks[19] ^ encoded_masks[20] ^ encoded_masks[26];
   assign decoded_masks_1[ 46] = encoded_masks[16] ^ encoded_masks[20] ^ encoded_masks[24];
   assign decoded_masks_1[ 47] = encoded_masks[23] ^ encoded_masks[28] ^ encoded_masks[29];
   assign decoded_masks_1[ 48] = encoded_masks[18] ^ encoded_masks[22] ^ encoded_masks[27];
   assign decoded_masks_1[ 49] = encoded_masks[15] ^ encoded_masks[19] ^ encoded_masks[25];
   assign decoded_masks_1[ 50] = encoded_masks[18] ^ encoded_masks[21] ^ encoded_masks[26];
   assign decoded_masks_1[ 51] = encoded_masks[17] ^ encoded_masks[19] ^ encoded_masks[27];
   assign decoded_masks_1[ 52] = encoded_masks[21] ^ encoded_masks[23] ^ encoded_masks[29];
   assign decoded_masks_1[ 53] = encoded_masks[17] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[ 54] = encoded_masks[22] ^ encoded_masks[26] ^ encoded_masks[29];
   assign decoded_masks_1[ 55] = encoded_masks[17] ^ encoded_masks[25] ^ encoded_masks[28];
   assign decoded_masks_1[ 56] = encoded_masks[16] ^ encoded_masks[20] ^ encoded_masks[27];
   assign decoded_masks_1[ 57] = encoded_masks[18] ^ encoded_masks[19] ^ encoded_masks[20];
   assign decoded_masks_1[ 58] = encoded_masks[23] ^ encoded_masks[24] ^ encoded_masks[25];
   assign decoded_masks_1[ 59] = encoded_masks[21] ^ encoded_masks[22] ^ encoded_masks[28];
   assign decoded_masks_1[ 60] = encoded_masks[20] ^ encoded_masks[22] ^ encoded_masks[25];
   assign decoded_masks_1[ 61] = encoded_masks[17] ^ encoded_masks[21] ^ encoded_masks[23];
   assign decoded_masks_1[ 62] = encoded_masks[15] ^ encoded_masks[24] ^ encoded_masks[28];
   assign decoded_masks_1[ 63] = encoded_masks[26] ^ encoded_masks[27] ^ encoded_masks[29];
   assign decoded_masks_1[ 64] = encoded_masks[18] ^ encoded_masks[20] ^ encoded_masks[23];
   assign decoded_masks_1[ 65] = encoded_masks[18] ^ encoded_masks[19] ^ encoded_masks[22];
   assign decoded_masks_1[ 66] = encoded_masks[15] ^ encoded_masks[24] ^ encoded_masks[29];
   assign decoded_masks_1[ 67] = encoded_masks[19] ^ encoded_masks[21] ^ encoded_masks[25];
   assign decoded_masks_1[ 68] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[28];
   assign decoded_masks_1[ 69] = encoded_masks[20] ^ encoded_masks[21] ^ encoded_masks[27];
   assign decoded_masks_1[ 70] = encoded_masks[17] ^ encoded_masks[23] ^ encoded_masks[26];
   assign decoded_masks_1[ 71] = encoded_masks[19] ^ encoded_masks[27] ^ encoded_masks[29];
   assign decoded_masks_1[ 72] = encoded_masks[15] ^ encoded_masks[18] ^ encoded_masks[22];
   assign decoded_masks_1[ 73] = encoded_masks[20] ^ encoded_masks[24] ^ encoded_masks[25];
   assign decoded_masks_1[ 74] = encoded_masks[15] ^ encoded_masks[21] ^ encoded_masks[26];
   assign decoded_masks_1[ 75] = encoded_masks[18] ^ encoded_masks[26] ^ encoded_masks[28];
   assign decoded_masks_1[ 76] = encoded_masks[22] ^ encoded_masks[24] ^ encoded_masks[27];
   assign decoded_masks_1[ 77] = encoded_masks[19] ^ encoded_masks[25] ^ encoded_masks[29];
   assign decoded_masks_1[ 78] = encoded_masks[18] ^ encoded_masks[23] ^ encoded_masks[24];
   assign decoded_masks_1[ 79] = encoded_masks[25] ^ encoded_masks[28] ^ encoded_masks[29];
   assign decoded_masks_1[ 80] = encoded_masks[17] ^ encoded_masks[20] ^ encoded_masks[21];
   assign decoded_masks_1[ 81] = encoded_masks[16] ^ encoded_masks[22] ^ encoded_masks[23];
   assign decoded_masks_1[ 82] = encoded_masks[20] ^ encoded_masks[26] ^ encoded_masks[27];
   assign decoded_masks_1[ 83] = encoded_masks[15] ^ encoded_masks[19] ^ encoded_masks[26];
   assign decoded_masks_1[ 84] = encoded_masks[17] ^ encoded_masks[19] ^ encoded_masks[22];
   assign decoded_masks_1[ 85] = encoded_masks[24] ^ encoded_masks[28] ^ encoded_masks[29];
   assign decoded_masks_1[ 86] = encoded_masks[16] ^ encoded_masks[21] ^ encoded_masks[25];
   assign decoded_masks_1[ 87] = encoded_masks[17] ^ encoded_masks[18] ^ encoded_masks[27];
   assign decoded_masks_1[ 88] = encoded_masks[19] ^ encoded_masks[24] ^ encoded_masks[28];
   assign decoded_masks_1[ 89] = encoded_masks[18] ^ encoded_masks[25] ^ encoded_masks[27];
   assign decoded_masks_1[ 90] = encoded_masks[20] ^ encoded_masks[23] ^ encoded_masks[28];
   assign decoded_masks_1[ 91] = encoded_masks[22] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[ 92] = encoded_masks[19] ^ encoded_masks[21] ^ encoded_masks[23];
   assign decoded_masks_1[ 93] = encoded_masks[15] ^ encoded_masks[17] ^ encoded_masks[29];
   assign decoded_masks_1[ 94] = encoded_masks[16] ^ encoded_masks[21] ^ encoded_masks[28];
   assign decoded_masks_1[ 95] = encoded_masks[23] ^ encoded_masks[25] ^ encoded_masks[29];
   assign decoded_masks_1[ 96] = encoded_masks[20] ^ encoded_masks[22] ^ encoded_masks[26];
   assign decoded_masks_1[ 97] = encoded_masks[17] ^ encoded_masks[18] ^ encoded_masks[24];
   assign decoded_masks_1[ 98] = encoded_masks[15] ^ encoded_masks[20] ^ encoded_masks[27];
   assign decoded_masks_1[ 99] = encoded_masks[18] ^ encoded_masks[23] ^ encoded_masks[25];
   assign decoded_masks_1[100] = encoded_masks[27] ^ encoded_masks[28] ^ encoded_masks[29];
   assign decoded_masks_1[101] = encoded_masks[19] ^ encoded_masks[20] ^ encoded_masks[22];
   assign decoded_masks_1[102] = encoded_masks[17] ^ encoded_masks[26] ^ encoded_masks[27];
   assign decoded_masks_1[103] = encoded_masks[16] ^ encoded_masks[19] ^ encoded_masks[25];
   assign decoded_masks_1[104] = encoded_masks[17] ^ encoded_masks[21] ^ encoded_masks[24];
   assign decoded_masks_1[105] = encoded_masks[22] ^ encoded_masks[25] ^ encoded_masks[26];
   assign decoded_masks_1[106] = encoded_masks[15] ^ encoded_masks[21] ^ encoded_masks[28];
   assign decoded_masks_1[107] = encoded_masks[18] ^ encoded_masks[19] ^ encoded_masks[29];
   assign decoded_masks_1[108] = encoded_masks[23] ^ encoded_masks[27] ^ encoded_masks[28];
   assign decoded_masks_1[109] = encoded_masks[16] ^ encoded_masks[22] ^ encoded_masks[26];
   assign decoded_masks_1[110] = encoded_masks[20] ^ encoded_masks[27] ^ encoded_masks[29];
   assign decoded_masks_1[111] = encoded_masks[20] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[112] = encoded_masks[15] ^ encoded_masks[22] ^ encoded_masks[23];
   assign decoded_masks_1[113] = encoded_masks[17] ^ encoded_masks[21] ^ encoded_masks[29];
   assign decoded_masks_1[114] = encoded_masks[17] ^ encoded_masks[18] ^ encoded_masks[28];
   assign decoded_masks_1[115] = encoded_masks[18] ^ encoded_masks[19] ^ encoded_masks[25];
   assign decoded_masks_1[116] = encoded_masks[15] ^ encoded_masks[23] ^ encoded_masks[26];
   assign decoded_masks_1[117] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[29];
   assign decoded_masks_1[118] = encoded_masks[21] ^ encoded_masks[23] ^ encoded_masks[27];
   assign decoded_masks_1[119] = encoded_masks[19] ^ encoded_masks[20] ^ encoded_masks[28];
   assign decoded_masks_1[120] = encoded_masks[17] ^ encoded_masks[24] ^ encoded_masks[25];
   assign decoded_masks_1[121] = encoded_masks[18] ^ encoded_masks[21] ^ encoded_masks[29];
   assign decoded_masks_1[122] = encoded_masks[19] ^ encoded_masks[23] ^ encoded_masks[24];
   assign decoded_masks_1[123] = encoded_masks[15] ^ encoded_masks[22] ^ encoded_masks[25];
   assign decoded_masks_1[124] = encoded_masks[18] ^ encoded_masks[21] ^ encoded_masks[27];
   assign decoded_masks_1[125] = encoded_masks[22] ^ encoded_masks[23] ^ encoded_masks[28];
   assign decoded_masks_1[126] = encoded_masks[16] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[127] = encoded_masks[20] ^ encoded_masks[26] ^ encoded_masks[28];
   assign decoded_masks_1[128] = encoded_masks[17] ^ encoded_masks[22] ^ encoded_masks[29];
   assign decoded_masks_1[129] = encoded_masks[16] ^ encoded_masks[18] ^ encoded_masks[25];
   assign decoded_masks_1[130] = encoded_masks[16] ^ encoded_masks[18] ^ encoded_masks[19];
   assign decoded_masks_1[131] = encoded_masks[21] ^ encoded_masks[24] ^ encoded_masks[26];
   assign decoded_masks_1[132] = encoded_masks[17] ^ encoded_masks[23] ^ encoded_masks[27];
   assign decoded_masks_1[133] = encoded_masks[15] ^ encoded_masks[20] ^ encoded_masks[28];
   assign decoded_masks_1[134] = encoded_masks[19] ^ encoded_masks[24] ^ encoded_masks[29];
   assign decoded_masks_1[135] = encoded_masks[15] ^ encoded_masks[20] ^ encoded_masks[21];
   assign decoded_masks_1[136] = encoded_masks[22] ^ encoded_masks[23] ^ encoded_masks[25];
   assign decoded_masks_1[137] = encoded_masks[25] ^ encoded_masks[27] ^ encoded_masks[28];
   assign decoded_masks_1[138] = encoded_masks[19] ^ encoded_masks[21] ^ encoded_masks[29];
   assign decoded_masks_1[139] = encoded_masks[16] ^ encoded_masks[22] ^ encoded_masks[24];
   assign decoded_masks_1[140] = encoded_masks[20] ^ encoded_masks[28] ^ encoded_masks[29];
   assign decoded_masks_1[141] = encoded_masks[19] ^ encoded_masks[26] ^ encoded_masks[27];
   assign decoded_masks_1[142] = encoded_masks[16] ^ encoded_masks[18] ^ encoded_masks[27];
   assign decoded_masks_1[143] = encoded_masks[17] ^ encoded_masks[18] ^ encoded_masks[26];
   assign decoded_masks_1[144] = encoded_masks[17] ^ encoded_masks[20] ^ encoded_masks[22];
   assign decoded_masks_1[145] = encoded_masks[15] ^ encoded_masks[21] ^ encoded_masks[25];
   assign decoded_masks_1[146] = encoded_masks[20] ^ encoded_masks[23] ^ encoded_masks[29];
   assign decoded_masks_1[147] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[24];
   assign decoded_masks_1[148] = encoded_masks[18] ^ encoded_masks[21] ^ encoded_masks[28];
   assign decoded_masks_1[149] = encoded_masks[22] ^ encoded_masks[23] ^ encoded_masks[24];
   assign decoded_masks_1[150] = encoded_masks[22] ^ encoded_masks[26] ^ encoded_masks[28];
   assign decoded_masks_1[151] = encoded_masks[20] ^ encoded_masks[26] ^ encoded_masks[29];
   assign decoded_masks_1[152] = encoded_masks[19] ^ encoded_masks[25] ^ encoded_masks[27];
   assign decoded_masks_1[153] = encoded_masks[15] ^ encoded_masks[18] ^ encoded_masks[23];
   assign decoded_masks_1[154] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[19];
   assign decoded_masks_1[155] = encoded_masks[21] ^ encoded_masks[24] ^ encoded_masks[27];
   assign decoded_masks_1[156] = encoded_masks[18] ^ encoded_masks[22] ^ encoded_masks[29];
   assign decoded_masks_1[157] = encoded_masks[22] ^ encoded_masks[24] ^ encoded_masks[25];
   assign decoded_masks_1[158] = encoded_masks[19] ^ encoded_masks[20] ^ encoded_masks[23];
   assign decoded_masks_1[159] = encoded_masks[15] ^ encoded_masks[26] ^ encoded_masks[27];
   assign decoded_masks_1[160] = encoded_masks[16] ^ encoded_masks[21] ^ encoded_masks[27];
   assign decoded_masks_1[161] = encoded_masks[25] ^ encoded_masks[26] ^ encoded_masks[28];
   assign decoded_masks_1[162] = encoded_masks[17] ^ encoded_masks[18] ^ encoded_masks[19];
   assign decoded_masks_1[163] = encoded_masks[21] ^ encoded_masks[24] ^ encoded_masks[28];
   assign decoded_masks_1[164] = encoded_masks[16] ^ encoded_masks[17] ^ encoded_masks[23];
   assign decoded_masks_1[165] = encoded_masks[17] ^ encoded_masks[20] ^ encoded_masks[25];
   assign decoded_masks_1[166] = encoded_masks[20] ^ encoded_masks[25] ^ encoded_masks[26];
   assign decoded_masks_1[167] = encoded_masks[18] ^ encoded_masks[24] ^ encoded_masks[29];
   assign decoded_masks_1[168] = encoded_masks[19] ^ encoded_masks[23] ^ encoded_masks[26];
   assign decoded_masks_1[169] = encoded_masks[22] ^ encoded_masks[25] ^ encoded_masks[27];
   assign decoded_masks_1[170] = encoded_masks[21] ^ encoded_masks[27] ^ encoded_masks[29];
   assign decoded_masks_1[171] = encoded_masks[15] ^ encoded_masks[19] ^ encoded_masks[24];
   assign decoded_masks_1[172] = encoded_masks[17] ^ encoded_masks[20] ^ encoded_masks[27];
   assign decoded_masks_1[173] = encoded_masks[16] ^ encoded_masks[21] ^ encoded_masks[22];
   assign decoded_masks_1[174] = encoded_masks[16] ^ encoded_masks[23] ^ encoded_masks[29];
   assign decoded_masks_1[175] = encoded_masks[15] ^ encoded_masks[17] ^ encoded_masks[28];
   assign decoded_masks_1[176] = encoded_masks[18] ^ encoded_masks[20] ^ encoded_masks[24];
   assign decoded_masks_1[177] = encoded_masks[15] ^ encoded_masks[19] ^ encoded_masks[28];
   assign decoded_masks_1[178] = encoded_masks[16] ^ encoded_masks[22] ^ encoded_masks[27];
   assign decoded_masks_1[179] = encoded_masks[15] ^ encoded_masks[18] ^ encoded_masks[29];
   assign decoded_masks_1[180] = encoded_masks[21] ^ encoded_masks[23] ^ encoded_masks[28];
   assign decoded_masks_1[181] = encoded_masks[17] ^ encoded_masks[21] ^ encoded_masks[25];
   assign decoded_masks_1[182] = encoded_masks[17] ^ encoded_masks[19] ^ encoded_masks[26];
   assign decoded_masks_1[183] = encoded_masks[20] ^ encoded_masks[24] ^ encoded_masks[28];
   assign decoded_masks_1[184] = encoded_masks[23] ^ encoded_masks[25] ^ encoded_masks[26];

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_controller (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire         edt_low_power_shift_en,
   input  wire [  3:0] edt_channels_in,
   input  wire [370:0] edt_decompressor_out,
   output wire [  3:0] edt_channels_out_from_controller,
   output wire [185:0] masks_for_compactor_0,
   output wire [184:0] masks_for_compactor_1,
   output wire [370:0] edt_scan_in
);
   reg    [  7:0] masks_shift_reg_0;
   reg    [  7:0] masks_shift_reg_1;
   reg    [  7:0] masks_shift_reg_2;
   reg    [  6:0] masks_shift_reg_3;
   reg    [  7:0] masks_hold_reg_0;
   reg    [  7:0] masks_hold_reg_1;
   reg    [  7:0] masks_hold_reg_2;
   reg    [  6:0] masks_hold_reg_3;
   wire           control_bit;
   wire   [  7:0] onehot_encoded_masks_0;
   wire   [  7:0] onehot_encoded_masks_1;
   wire   [ 29:0] xor_encoded_masks;
   wire   [185:0] onehot_decoded_masks_0;
   wire   [184:0] onehot_decoded_masks_1;
   wire   [185:0] xor_decoded_masks_0;
   wire   [184:0] xor_decoded_masks_1;
   wire           masks_shift_reg_sync_reset;
   wire   [  3:0] edt_channels_out_from_low_power_shift_control;

   firebird7_in_gate2_tessent_edt_intest_edt_low_power_shift_controller low_power_shift_controller_i (
      .edt_clock(edt_clock),
      .edt_update(edt_update),
      .edt_low_power_shift_en(edt_low_power_shift_en),
      .edt_channels_in(edt_channels_in),
      .edt_decompressor_out(edt_decompressor_out),
      .edt_channels_out_from_low_power_shift_control(edt_channels_out_from_low_power_shift_control),
      .edt_scan_in(edt_scan_in));

   assign masks_shift_reg_sync_reset = edt_update;

   // synopsys sync_set_reset masks_shift_reg_sync_reset
   always @(posedge edt_clock)
   begin : shift_masks_regs
      if (masks_shift_reg_sync_reset == 1'b1) begin
         masks_shift_reg_0 <= 8'b00000000;
         masks_shift_reg_1 <= 8'b00000000;
         masks_shift_reg_2 <= 8'b00000000;
         masks_shift_reg_3 <= 7'b0000000;
      end
      else begin
         masks_shift_reg_0 <= {edt_channels_out_from_low_power_shift_control[0], masks_shift_reg_0[7:1]};
         masks_shift_reg_1 <= {edt_channels_out_from_low_power_shift_control[1], masks_shift_reg_1[7:1]};
         masks_shift_reg_2 <= {edt_channels_out_from_low_power_shift_control[2], masks_shift_reg_2[7:1]};
         masks_shift_reg_3 <= {edt_channels_out_from_low_power_shift_control[3], masks_shift_reg_3[6:1]};
      end
   end

   always @(posedge edt_clock)
   begin : update_masks_regs
      if (edt_update == 1'b1) begin
         masks_hold_reg_0 <= masks_shift_reg_0;
         masks_hold_reg_1 <= masks_shift_reg_1;
         masks_hold_reg_2 <= masks_shift_reg_2;
         masks_hold_reg_3 <= masks_shift_reg_3;
      end
   end

   assign edt_channels_out_from_controller[0] = masks_shift_reg_0[0];
   assign edt_channels_out_from_controller[1] = masks_shift_reg_1[0];
   assign edt_channels_out_from_controller[2] = masks_shift_reg_2[0];
   assign edt_channels_out_from_controller[3] = masks_shift_reg_3[0];

   assign control_bit = masks_hold_reg_0[7];

   assign xor_encoded_masks = {masks_hold_reg_3[0], masks_hold_reg_3[1], masks_hold_reg_3[2], 
                               masks_hold_reg_3[3], masks_hold_reg_3[4], masks_hold_reg_3[5], 
                               masks_hold_reg_3[6], masks_hold_reg_2[0], masks_hold_reg_2[1], 
                               masks_hold_reg_2[2], masks_hold_reg_2[3], masks_hold_reg_2[4], 
                               masks_hold_reg_2[5], masks_hold_reg_2[6], masks_hold_reg_2[7], 
                               masks_hold_reg_1[0], masks_hold_reg_1[1], masks_hold_reg_1[2], 
                               masks_hold_reg_1[3], masks_hold_reg_1[4], masks_hold_reg_1[5], 
                               masks_hold_reg_1[6], masks_hold_reg_1[7], masks_hold_reg_0[0], 
                               masks_hold_reg_0[1], masks_hold_reg_0[2], masks_hold_reg_0[3], 
                               masks_hold_reg_0[4], masks_hold_reg_0[5], masks_hold_reg_0[6]};

   assign onehot_encoded_masks_0 = {masks_hold_reg_0[6], masks_hold_reg_0[5], masks_hold_reg_0[4], 
                                    masks_hold_reg_0[3], masks_hold_reg_0[2], masks_hold_reg_0[1], 
                                    masks_hold_reg_0[0], masks_hold_reg_1[7]};
   assign onehot_encoded_masks_1 = {masks_hold_reg_2[7], masks_hold_reg_2[6], masks_hold_reg_2[5], 
                                    masks_hold_reg_2[4], masks_hold_reg_2[3], masks_hold_reg_2[2], 
                                    masks_hold_reg_2[1], masks_hold_reg_2[0]};

   firebird7_in_gate2_tessent_edt_intest_edt_xor_decoder xor_decoder (
      .encoded_masks(xor_encoded_masks),
      .decoded_masks_0(xor_decoded_masks_0),
      .decoded_masks_1(xor_decoded_masks_1));

   firebird7_in_gate2_tessent_edt_intest_edt_onehot_decoder_8_to_186 decoder1 (.encoded_masks(onehot_encoded_masks_0),
                                                                               .decoded_masks(onehot_decoded_masks_0));
   firebird7_in_gate2_tessent_edt_intest_edt_onehot_decoder_8_to_185 decoder2 (.encoded_masks(onehot_encoded_masks_1),
                                                                               .decoded_masks(onehot_decoded_masks_1));

   assign masks_for_compactor_0 = control_bit ? onehot_decoded_masks_0 : xor_decoded_masks_0;
   assign masks_for_compactor_1 = control_bit ? onehot_decoded_masks_1 : xor_decoded_masks_1;
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_spatial_compactor_185_w_output_lockup (
   input  wire         edt_clock,
   input  wire [184:0] multi_bit_input,
   output reg          single_bit_output
);
   reg    [ 92:0] level1;
   reg    [ 46:0] level2;
   reg    [ 23:0] level3;
   reg    [ 11:0] level4;
   reg    [  5:0] level5;
   reg    [  2:0] level6;
   reg    [  1:0] level7;
   reg            level8_pipelined;

   always @(multi_bit_input)
   begin : compact185_level1
      level1[ 0] = multi_bit_input[  0] ^ multi_bit_input[  1];
      level1[ 1] = multi_bit_input[  2] ^ multi_bit_input[  3];
      level1[ 2] = multi_bit_input[  4] ^ multi_bit_input[  5];
      level1[ 3] = multi_bit_input[  6] ^ multi_bit_input[  7];
      level1[ 4] = multi_bit_input[  8] ^ multi_bit_input[  9];
      level1[ 5] = multi_bit_input[ 10] ^ multi_bit_input[ 11];
      level1[ 6] = multi_bit_input[ 12] ^ multi_bit_input[ 13];
      level1[ 7] = multi_bit_input[ 14] ^ multi_bit_input[ 15];
      level1[ 8] = multi_bit_input[ 16] ^ multi_bit_input[ 17];
      level1[ 9] = multi_bit_input[ 18] ^ multi_bit_input[ 19];
      level1[10] = multi_bit_input[ 20] ^ multi_bit_input[ 21];
      level1[11] = multi_bit_input[ 22] ^ multi_bit_input[ 23];
      level1[12] = multi_bit_input[ 24] ^ multi_bit_input[ 25];
      level1[13] = multi_bit_input[ 26] ^ multi_bit_input[ 27];
      level1[14] = multi_bit_input[ 28] ^ multi_bit_input[ 29];
      level1[15] = multi_bit_input[ 30] ^ multi_bit_input[ 31];
      level1[16] = multi_bit_input[ 32] ^ multi_bit_input[ 33];
      level1[17] = multi_bit_input[ 34] ^ multi_bit_input[ 35];
      level1[18] = multi_bit_input[ 36] ^ multi_bit_input[ 37];
      level1[19] = multi_bit_input[ 38] ^ multi_bit_input[ 39];
      level1[20] = multi_bit_input[ 40] ^ multi_bit_input[ 41];
      level1[21] = multi_bit_input[ 42] ^ multi_bit_input[ 43];
      level1[22] = multi_bit_input[ 44] ^ multi_bit_input[ 45];
      level1[23] = multi_bit_input[ 46] ^ multi_bit_input[ 47];
      level1[24] = multi_bit_input[ 48] ^ multi_bit_input[ 49];
      level1[25] = multi_bit_input[ 50] ^ multi_bit_input[ 51];
      level1[26] = multi_bit_input[ 52] ^ multi_bit_input[ 53];
      level1[27] = multi_bit_input[ 54] ^ multi_bit_input[ 55];
      level1[28] = multi_bit_input[ 56] ^ multi_bit_input[ 57];
      level1[29] = multi_bit_input[ 58] ^ multi_bit_input[ 59];
      level1[30] = multi_bit_input[ 60] ^ multi_bit_input[ 61];
      level1[31] = multi_bit_input[ 62] ^ multi_bit_input[ 63];
      level1[32] = multi_bit_input[ 64] ^ multi_bit_input[ 65];
      level1[33] = multi_bit_input[ 66] ^ multi_bit_input[ 67];
      level1[34] = multi_bit_input[ 68] ^ multi_bit_input[ 69];
      level1[35] = multi_bit_input[ 70] ^ multi_bit_input[ 71];
      level1[36] = multi_bit_input[ 72] ^ multi_bit_input[ 73];
      level1[37] = multi_bit_input[ 74] ^ multi_bit_input[ 75];
      level1[38] = multi_bit_input[ 76] ^ multi_bit_input[ 77];
      level1[39] = multi_bit_input[ 78] ^ multi_bit_input[ 79];
      level1[40] = multi_bit_input[ 80] ^ multi_bit_input[ 81];
      level1[41] = multi_bit_input[ 82] ^ multi_bit_input[ 83];
      level1[42] = multi_bit_input[ 84] ^ multi_bit_input[ 85];
      level1[43] = multi_bit_input[ 86] ^ multi_bit_input[ 87];
      level1[44] = multi_bit_input[ 88] ^ multi_bit_input[ 89];
      level1[45] = multi_bit_input[ 90] ^ multi_bit_input[ 91];
      level1[46] = multi_bit_input[ 92] ^ multi_bit_input[ 93];
      level1[47] = multi_bit_input[ 94] ^ multi_bit_input[ 95];
      level1[48] = multi_bit_input[ 96] ^ multi_bit_input[ 97];
      level1[49] = multi_bit_input[ 98] ^ multi_bit_input[ 99];
      level1[50] = multi_bit_input[100] ^ multi_bit_input[101];
      level1[51] = multi_bit_input[102] ^ multi_bit_input[103];
      level1[52] = multi_bit_input[104] ^ multi_bit_input[105];
      level1[53] = multi_bit_input[106] ^ multi_bit_input[107];
      level1[54] = multi_bit_input[108] ^ multi_bit_input[109];
      level1[55] = multi_bit_input[110] ^ multi_bit_input[111];
      level1[56] = multi_bit_input[112] ^ multi_bit_input[113];
      level1[57] = multi_bit_input[114] ^ multi_bit_input[115];
      level1[58] = multi_bit_input[116] ^ multi_bit_input[117];
      level1[59] = multi_bit_input[118] ^ multi_bit_input[119];
      level1[60] = multi_bit_input[120] ^ multi_bit_input[121];
      level1[61] = multi_bit_input[122] ^ multi_bit_input[123];
      level1[62] = multi_bit_input[124] ^ multi_bit_input[125];
      level1[63] = multi_bit_input[126] ^ multi_bit_input[127];
      level1[64] = multi_bit_input[128] ^ multi_bit_input[129];
      level1[65] = multi_bit_input[130] ^ multi_bit_input[131];
      level1[66] = multi_bit_input[132] ^ multi_bit_input[133];
      level1[67] = multi_bit_input[134] ^ multi_bit_input[135];
      level1[68] = multi_bit_input[136] ^ multi_bit_input[137];
      level1[69] = multi_bit_input[138] ^ multi_bit_input[139];
      level1[70] = multi_bit_input[140] ^ multi_bit_input[141];
      level1[71] = multi_bit_input[142] ^ multi_bit_input[143];
      level1[72] = multi_bit_input[144] ^ multi_bit_input[145];
      level1[73] = multi_bit_input[146] ^ multi_bit_input[147];
      level1[74] = multi_bit_input[148] ^ multi_bit_input[149];
      level1[75] = multi_bit_input[150] ^ multi_bit_input[151];
      level1[76] = multi_bit_input[152] ^ multi_bit_input[153];
      level1[77] = multi_bit_input[154] ^ multi_bit_input[155];
      level1[78] = multi_bit_input[156] ^ multi_bit_input[157];
      level1[79] = multi_bit_input[158] ^ multi_bit_input[159];
      level1[80] = multi_bit_input[160] ^ multi_bit_input[161];
      level1[81] = multi_bit_input[162] ^ multi_bit_input[163];
      level1[82] = multi_bit_input[164] ^ multi_bit_input[165];
      level1[83] = multi_bit_input[166] ^ multi_bit_input[167];
      level1[84] = multi_bit_input[168] ^ multi_bit_input[169];
      level1[85] = multi_bit_input[170] ^ multi_bit_input[171];
      level1[86] = multi_bit_input[172] ^ multi_bit_input[173];
      level1[87] = multi_bit_input[174] ^ multi_bit_input[175];
      level1[88] = multi_bit_input[176] ^ multi_bit_input[177];
      level1[89] = multi_bit_input[178] ^ multi_bit_input[179];
      level1[90] = multi_bit_input[180] ^ multi_bit_input[181];
      level1[91] = multi_bit_input[182] ^ multi_bit_input[183];
      level1[92] = multi_bit_input[184];
   end

   always @(level1)
   begin : compact185_level2
      level2[ 0] = level1[ 0] ^ level1[ 1];
      level2[ 1] = level1[ 2] ^ level1[ 3];
      level2[ 2] = level1[ 4] ^ level1[ 5];
      level2[ 3] = level1[ 6] ^ level1[ 7];
      level2[ 4] = level1[ 8] ^ level1[ 9];
      level2[ 5] = level1[10] ^ level1[11];
      level2[ 6] = level1[12] ^ level1[13];
      level2[ 7] = level1[14] ^ level1[15];
      level2[ 8] = level1[16] ^ level1[17];
      level2[ 9] = level1[18] ^ level1[19];
      level2[10] = level1[20] ^ level1[21];
      level2[11] = level1[22] ^ level1[23];
      level2[12] = level1[24] ^ level1[25];
      level2[13] = level1[26] ^ level1[27];
      level2[14] = level1[28] ^ level1[29];
      level2[15] = level1[30] ^ level1[31];
      level2[16] = level1[32] ^ level1[33];
      level2[17] = level1[34] ^ level1[35];
      level2[18] = level1[36] ^ level1[37];
      level2[19] = level1[38] ^ level1[39];
      level2[20] = level1[40] ^ level1[41];
      level2[21] = level1[42] ^ level1[43];
      level2[22] = level1[44] ^ level1[45];
      level2[23] = level1[46] ^ level1[47];
      level2[24] = level1[48] ^ level1[49];
      level2[25] = level1[50] ^ level1[51];
      level2[26] = level1[52] ^ level1[53];
      level2[27] = level1[54] ^ level1[55];
      level2[28] = level1[56] ^ level1[57];
      level2[29] = level1[58] ^ level1[59];
      level2[30] = level1[60] ^ level1[61];
      level2[31] = level1[62] ^ level1[63];
      level2[32] = level1[64] ^ level1[65];
      level2[33] = level1[66] ^ level1[67];
      level2[34] = level1[68] ^ level1[69];
      level2[35] = level1[70] ^ level1[71];
      level2[36] = level1[72] ^ level1[73];
      level2[37] = level1[74] ^ level1[75];
      level2[38] = level1[76] ^ level1[77];
      level2[39] = level1[78] ^ level1[79];
      level2[40] = level1[80] ^ level1[81];
      level2[41] = level1[82] ^ level1[83];
      level2[42] = level1[84] ^ level1[85];
      level2[43] = level1[86] ^ level1[87];
      level2[44] = level1[88] ^ level1[89];
      level2[45] = level1[90] ^ level1[91];
      level2[46] = level1[92];
   end

   always @(level2)
   begin : compact185_level3
      level3[ 0] = level2[ 0] ^ level2[ 1];
      level3[ 1] = level2[ 2] ^ level2[ 3];
      level3[ 2] = level2[ 4] ^ level2[ 5];
      level3[ 3] = level2[ 6] ^ level2[ 7];
      level3[ 4] = level2[ 8] ^ level2[ 9];
      level3[ 5] = level2[10] ^ level2[11];
      level3[ 6] = level2[12] ^ level2[13];
      level3[ 7] = level2[14] ^ level2[15];
      level3[ 8] = level2[16] ^ level2[17];
      level3[ 9] = level2[18] ^ level2[19];
      level3[10] = level2[20] ^ level2[21];
      level3[11] = level2[22] ^ level2[23];
      level3[12] = level2[24] ^ level2[25];
      level3[13] = level2[26] ^ level2[27];
      level3[14] = level2[28] ^ level2[29];
      level3[15] = level2[30] ^ level2[31];
      level3[16] = level2[32] ^ level2[33];
      level3[17] = level2[34] ^ level2[35];
      level3[18] = level2[36] ^ level2[37];
      level3[19] = level2[38] ^ level2[39];
      level3[20] = level2[40] ^ level2[41];
      level3[21] = level2[42] ^ level2[43];
      level3[22] = level2[44] ^ level2[45];
      level3[23] = level2[46];
   end

   always @(level3)
   begin : compact185_level4
      level4[ 0] = level3[ 0] ^ level3[ 1];
      level4[ 1] = level3[ 2] ^ level3[ 3];
      level4[ 2] = level3[ 4] ^ level3[ 5];
      level4[ 3] = level3[ 6] ^ level3[ 7];
      level4[ 4] = level3[ 8] ^ level3[ 9];
      level4[ 5] = level3[10] ^ level3[11];
      level4[ 6] = level3[12] ^ level3[13];
      level4[ 7] = level3[14] ^ level3[15];
      level4[ 8] = level3[16] ^ level3[17];
      level4[ 9] = level3[18] ^ level3[19];
      level4[10] = level3[20] ^ level3[21];
      level4[11] = level3[22] ^ level3[23];
   end

   always @(level4)
   begin : compact185_level5
      level5[0] = level4[ 0] ^ level4[ 1];
      level5[1] = level4[ 2] ^ level4[ 3];
      level5[2] = level4[ 4] ^ level4[ 5];
      level5[3] = level4[ 6] ^ level4[ 7];
      level5[4] = level4[ 8] ^ level4[ 9];
      level5[5] = level4[10] ^ level4[11];
   end

   always @(level5)
   begin : compact185_level6
      level6[0] = level5[0] ^ level5[1];
      level6[1] = level5[2] ^ level5[3];
      level6[2] = level5[4] ^ level5[5];
   end

   always @(level6)
   begin : compact185_level7
      level7[0] = level6[0] ^ level6[1];
      level7[1] = level6[2];
   end

   always @(posedge edt_clock)
   begin : compact185_level8_pipelined
      level8_pipelined <= level7[0] ^ level7[1];
   end

   always @(negedge edt_clock)
   begin : compact185_level8_lockup
      single_bit_output <= level8_pipelined;
   end

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_spatial_compactor_186_w_output_lockup (
   input  wire         edt_clock,
   input  wire [185:0] multi_bit_input,
   output reg          single_bit_output
);
   reg    [ 92:0] level1;
   reg    [ 46:0] level2;
   reg    [ 23:0] level3;
   reg    [ 11:0] level4;
   reg    [  5:0] level5;
   reg    [  2:0] level6;
   reg    [  1:0] level7;
   reg            level8_pipelined;

   always @(multi_bit_input)
   begin : compact186_level1
      level1[ 0] = multi_bit_input[  0] ^ multi_bit_input[  1];
      level1[ 1] = multi_bit_input[  2] ^ multi_bit_input[  3];
      level1[ 2] = multi_bit_input[  4] ^ multi_bit_input[  5];
      level1[ 3] = multi_bit_input[  6] ^ multi_bit_input[  7];
      level1[ 4] = multi_bit_input[  8] ^ multi_bit_input[  9];
      level1[ 5] = multi_bit_input[ 10] ^ multi_bit_input[ 11];
      level1[ 6] = multi_bit_input[ 12] ^ multi_bit_input[ 13];
      level1[ 7] = multi_bit_input[ 14] ^ multi_bit_input[ 15];
      level1[ 8] = multi_bit_input[ 16] ^ multi_bit_input[ 17];
      level1[ 9] = multi_bit_input[ 18] ^ multi_bit_input[ 19];
      level1[10] = multi_bit_input[ 20] ^ multi_bit_input[ 21];
      level1[11] = multi_bit_input[ 22] ^ multi_bit_input[ 23];
      level1[12] = multi_bit_input[ 24] ^ multi_bit_input[ 25];
      level1[13] = multi_bit_input[ 26] ^ multi_bit_input[ 27];
      level1[14] = multi_bit_input[ 28] ^ multi_bit_input[ 29];
      level1[15] = multi_bit_input[ 30] ^ multi_bit_input[ 31];
      level1[16] = multi_bit_input[ 32] ^ multi_bit_input[ 33];
      level1[17] = multi_bit_input[ 34] ^ multi_bit_input[ 35];
      level1[18] = multi_bit_input[ 36] ^ multi_bit_input[ 37];
      level1[19] = multi_bit_input[ 38] ^ multi_bit_input[ 39];
      level1[20] = multi_bit_input[ 40] ^ multi_bit_input[ 41];
      level1[21] = multi_bit_input[ 42] ^ multi_bit_input[ 43];
      level1[22] = multi_bit_input[ 44] ^ multi_bit_input[ 45];
      level1[23] = multi_bit_input[ 46] ^ multi_bit_input[ 47];
      level1[24] = multi_bit_input[ 48] ^ multi_bit_input[ 49];
      level1[25] = multi_bit_input[ 50] ^ multi_bit_input[ 51];
      level1[26] = multi_bit_input[ 52] ^ multi_bit_input[ 53];
      level1[27] = multi_bit_input[ 54] ^ multi_bit_input[ 55];
      level1[28] = multi_bit_input[ 56] ^ multi_bit_input[ 57];
      level1[29] = multi_bit_input[ 58] ^ multi_bit_input[ 59];
      level1[30] = multi_bit_input[ 60] ^ multi_bit_input[ 61];
      level1[31] = multi_bit_input[ 62] ^ multi_bit_input[ 63];
      level1[32] = multi_bit_input[ 64] ^ multi_bit_input[ 65];
      level1[33] = multi_bit_input[ 66] ^ multi_bit_input[ 67];
      level1[34] = multi_bit_input[ 68] ^ multi_bit_input[ 69];
      level1[35] = multi_bit_input[ 70] ^ multi_bit_input[ 71];
      level1[36] = multi_bit_input[ 72] ^ multi_bit_input[ 73];
      level1[37] = multi_bit_input[ 74] ^ multi_bit_input[ 75];
      level1[38] = multi_bit_input[ 76] ^ multi_bit_input[ 77];
      level1[39] = multi_bit_input[ 78] ^ multi_bit_input[ 79];
      level1[40] = multi_bit_input[ 80] ^ multi_bit_input[ 81];
      level1[41] = multi_bit_input[ 82] ^ multi_bit_input[ 83];
      level1[42] = multi_bit_input[ 84] ^ multi_bit_input[ 85];
      level1[43] = multi_bit_input[ 86] ^ multi_bit_input[ 87];
      level1[44] = multi_bit_input[ 88] ^ multi_bit_input[ 89];
      level1[45] = multi_bit_input[ 90] ^ multi_bit_input[ 91];
      level1[46] = multi_bit_input[ 92] ^ multi_bit_input[ 93];
      level1[47] = multi_bit_input[ 94] ^ multi_bit_input[ 95];
      level1[48] = multi_bit_input[ 96] ^ multi_bit_input[ 97];
      level1[49] = multi_bit_input[ 98] ^ multi_bit_input[ 99];
      level1[50] = multi_bit_input[100] ^ multi_bit_input[101];
      level1[51] = multi_bit_input[102] ^ multi_bit_input[103];
      level1[52] = multi_bit_input[104] ^ multi_bit_input[105];
      level1[53] = multi_bit_input[106] ^ multi_bit_input[107];
      level1[54] = multi_bit_input[108] ^ multi_bit_input[109];
      level1[55] = multi_bit_input[110] ^ multi_bit_input[111];
      level1[56] = multi_bit_input[112] ^ multi_bit_input[113];
      level1[57] = multi_bit_input[114] ^ multi_bit_input[115];
      level1[58] = multi_bit_input[116] ^ multi_bit_input[117];
      level1[59] = multi_bit_input[118] ^ multi_bit_input[119];
      level1[60] = multi_bit_input[120] ^ multi_bit_input[121];
      level1[61] = multi_bit_input[122] ^ multi_bit_input[123];
      level1[62] = multi_bit_input[124] ^ multi_bit_input[125];
      level1[63] = multi_bit_input[126] ^ multi_bit_input[127];
      level1[64] = multi_bit_input[128] ^ multi_bit_input[129];
      level1[65] = multi_bit_input[130] ^ multi_bit_input[131];
      level1[66] = multi_bit_input[132] ^ multi_bit_input[133];
      level1[67] = multi_bit_input[134] ^ multi_bit_input[135];
      level1[68] = multi_bit_input[136] ^ multi_bit_input[137];
      level1[69] = multi_bit_input[138] ^ multi_bit_input[139];
      level1[70] = multi_bit_input[140] ^ multi_bit_input[141];
      level1[71] = multi_bit_input[142] ^ multi_bit_input[143];
      level1[72] = multi_bit_input[144] ^ multi_bit_input[145];
      level1[73] = multi_bit_input[146] ^ multi_bit_input[147];
      level1[74] = multi_bit_input[148] ^ multi_bit_input[149];
      level1[75] = multi_bit_input[150] ^ multi_bit_input[151];
      level1[76] = multi_bit_input[152] ^ multi_bit_input[153];
      level1[77] = multi_bit_input[154] ^ multi_bit_input[155];
      level1[78] = multi_bit_input[156] ^ multi_bit_input[157];
      level1[79] = multi_bit_input[158] ^ multi_bit_input[159];
      level1[80] = multi_bit_input[160] ^ multi_bit_input[161];
      level1[81] = multi_bit_input[162] ^ multi_bit_input[163];
      level1[82] = multi_bit_input[164] ^ multi_bit_input[165];
      level1[83] = multi_bit_input[166] ^ multi_bit_input[167];
      level1[84] = multi_bit_input[168] ^ multi_bit_input[169];
      level1[85] = multi_bit_input[170] ^ multi_bit_input[171];
      level1[86] = multi_bit_input[172] ^ multi_bit_input[173];
      level1[87] = multi_bit_input[174] ^ multi_bit_input[175];
      level1[88] = multi_bit_input[176] ^ multi_bit_input[177];
      level1[89] = multi_bit_input[178] ^ multi_bit_input[179];
      level1[90] = multi_bit_input[180] ^ multi_bit_input[181];
      level1[91] = multi_bit_input[182] ^ multi_bit_input[183];
      level1[92] = multi_bit_input[184] ^ multi_bit_input[185];
   end

   always @(level1)
   begin : compact186_level2
      level2[ 0] = level1[ 0] ^ level1[ 1];
      level2[ 1] = level1[ 2] ^ level1[ 3];
      level2[ 2] = level1[ 4] ^ level1[ 5];
      level2[ 3] = level1[ 6] ^ level1[ 7];
      level2[ 4] = level1[ 8] ^ level1[ 9];
      level2[ 5] = level1[10] ^ level1[11];
      level2[ 6] = level1[12] ^ level1[13];
      level2[ 7] = level1[14] ^ level1[15];
      level2[ 8] = level1[16] ^ level1[17];
      level2[ 9] = level1[18] ^ level1[19];
      level2[10] = level1[20] ^ level1[21];
      level2[11] = level1[22] ^ level1[23];
      level2[12] = level1[24] ^ level1[25];
      level2[13] = level1[26] ^ level1[27];
      level2[14] = level1[28] ^ level1[29];
      level2[15] = level1[30] ^ level1[31];
      level2[16] = level1[32] ^ level1[33];
      level2[17] = level1[34] ^ level1[35];
      level2[18] = level1[36] ^ level1[37];
      level2[19] = level1[38] ^ level1[39];
      level2[20] = level1[40] ^ level1[41];
      level2[21] = level1[42] ^ level1[43];
      level2[22] = level1[44] ^ level1[45];
      level2[23] = level1[46] ^ level1[47];
      level2[24] = level1[48] ^ level1[49];
      level2[25] = level1[50] ^ level1[51];
      level2[26] = level1[52] ^ level1[53];
      level2[27] = level1[54] ^ level1[55];
      level2[28] = level1[56] ^ level1[57];
      level2[29] = level1[58] ^ level1[59];
      level2[30] = level1[60] ^ level1[61];
      level2[31] = level1[62] ^ level1[63];
      level2[32] = level1[64] ^ level1[65];
      level2[33] = level1[66] ^ level1[67];
      level2[34] = level1[68] ^ level1[69];
      level2[35] = level1[70] ^ level1[71];
      level2[36] = level1[72] ^ level1[73];
      level2[37] = level1[74] ^ level1[75];
      level2[38] = level1[76] ^ level1[77];
      level2[39] = level1[78] ^ level1[79];
      level2[40] = level1[80] ^ level1[81];
      level2[41] = level1[82] ^ level1[83];
      level2[42] = level1[84] ^ level1[85];
      level2[43] = level1[86] ^ level1[87];
      level2[44] = level1[88] ^ level1[89];
      level2[45] = level1[90] ^ level1[91];
      level2[46] = level1[92];
   end

   always @(level2)
   begin : compact186_level3
      level3[ 0] = level2[ 0] ^ level2[ 1];
      level3[ 1] = level2[ 2] ^ level2[ 3];
      level3[ 2] = level2[ 4] ^ level2[ 5];
      level3[ 3] = level2[ 6] ^ level2[ 7];
      level3[ 4] = level2[ 8] ^ level2[ 9];
      level3[ 5] = level2[10] ^ level2[11];
      level3[ 6] = level2[12] ^ level2[13];
      level3[ 7] = level2[14] ^ level2[15];
      level3[ 8] = level2[16] ^ level2[17];
      level3[ 9] = level2[18] ^ level2[19];
      level3[10] = level2[20] ^ level2[21];
      level3[11] = level2[22] ^ level2[23];
      level3[12] = level2[24] ^ level2[25];
      level3[13] = level2[26] ^ level2[27];
      level3[14] = level2[28] ^ level2[29];
      level3[15] = level2[30] ^ level2[31];
      level3[16] = level2[32] ^ level2[33];
      level3[17] = level2[34] ^ level2[35];
      level3[18] = level2[36] ^ level2[37];
      level3[19] = level2[38] ^ level2[39];
      level3[20] = level2[40] ^ level2[41];
      level3[21] = level2[42] ^ level2[43];
      level3[22] = level2[44] ^ level2[45];
      level3[23] = level2[46];
   end

   always @(level3)
   begin : compact186_level4
      level4[ 0] = level3[ 0] ^ level3[ 1];
      level4[ 1] = level3[ 2] ^ level3[ 3];
      level4[ 2] = level3[ 4] ^ level3[ 5];
      level4[ 3] = level3[ 6] ^ level3[ 7];
      level4[ 4] = level3[ 8] ^ level3[ 9];
      level4[ 5] = level3[10] ^ level3[11];
      level4[ 6] = level3[12] ^ level3[13];
      level4[ 7] = level3[14] ^ level3[15];
      level4[ 8] = level3[16] ^ level3[17];
      level4[ 9] = level3[18] ^ level3[19];
      level4[10] = level3[20] ^ level3[21];
      level4[11] = level3[22] ^ level3[23];
   end

   always @(level4)
   begin : compact186_level5
      level5[0] = level4[ 0] ^ level4[ 1];
      level5[1] = level4[ 2] ^ level4[ 3];
      level5[2] = level4[ 4] ^ level4[ 5];
      level5[3] = level4[ 6] ^ level4[ 7];
      level5[4] = level4[ 8] ^ level4[ 9];
      level5[5] = level4[10] ^ level4[11];
   end

   always @(level5)
   begin : compact186_level6
      level6[0] = level5[0] ^ level5[1];
      level6[1] = level5[2] ^ level5[3];
      level6[2] = level5[4] ^ level5[5];
   end

   always @(level6)
   begin : compact186_level7
      level7[0] = level6[0] ^ level6[1];
      level7[1] = level6[2];
   end

   always @(posedge edt_clock)
   begin : compact186_level8_pipelined
      level8_pipelined <= level7[0] ^ level7[1];
   end

   always @(negedge edt_clock)
   begin : compact186_level8_lockup
      single_bit_output <= level8_pipelined;
   end

endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_compactor (
   input  wire         edt_clock,
   input  wire [370:0] edt_scan_out,
   input  wire [185:0] masks_for_compactor_0,
   input  wire [184:0] masks_for_compactor_1,
   output wire [  1:0] edt_channels_out
);
   wire   [185:0] masked_scan_outputs_0;
   wire   [184:0] masked_scan_outputs_1;

   assign masked_scan_outputs_0 = edt_scan_out[185:  0] & masks_for_compactor_0;
   assign masked_scan_outputs_1 = edt_scan_out[370:186] & masks_for_compactor_1;

   firebird7_in_gate2_tessent_edt_intest_edt_spatial_compactor_186_w_output_lockup compactor1 (.edt_clock(edt_clock),
                                                                                               .multi_bit_input(masked_scan_outputs_0),
                                                                                               .single_bit_output(edt_channels_out[0]));
   firebird7_in_gate2_tessent_edt_intest_edt_spatial_compactor_185_w_output_lockup compactor2 (.edt_clock(edt_clock),
                                                                                               .multi_bit_input(masked_scan_outputs_1),
                                                                                               .single_bit_output(edt_channels_out[1]));
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt_bypass_logic (
   input  wire         edt_bypass,
   input  wire [  3:0] edt_channels_in,
   output wire [  1:0] edt_channels_out,
   output wire [370:0] edt_scan_in,
   input  wire [370:0] edt_scan_out,
   input  wire [370:0] edt_bypass_in,
   input  wire [  1:0] edt_bypass_out
);

   assign edt_scan_in[0] = edt_bypass ? edt_channels_in[0] : edt_bypass_in[0];
   assign edt_scan_in[1] = edt_bypass ? edt_scan_out[0] : edt_bypass_in[1];
   assign edt_scan_in[2] = edt_bypass ? edt_scan_out[1] : edt_bypass_in[2];
   assign edt_scan_in[3] = edt_bypass ? edt_scan_out[2] : edt_bypass_in[3];
   assign edt_scan_in[4] = edt_bypass ? edt_scan_out[3] : edt_bypass_in[4];
   assign edt_scan_in[5] = edt_bypass ? edt_scan_out[4] : edt_bypass_in[5];
   assign edt_scan_in[6] = edt_bypass ? edt_scan_out[5] : edt_bypass_in[6];
   assign edt_scan_in[7] = edt_bypass ? edt_scan_out[6] : edt_bypass_in[7];
   assign edt_scan_in[8] = edt_bypass ? edt_scan_out[7] : edt_bypass_in[8];
   assign edt_scan_in[9] = edt_bypass ? edt_scan_out[8] : edt_bypass_in[9];
   assign edt_scan_in[10] = edt_bypass ? edt_scan_out[9] : edt_bypass_in[10];
   assign edt_scan_in[11] = edt_bypass ? edt_scan_out[10] : edt_bypass_in[11];
   assign edt_scan_in[12] = edt_bypass ? edt_scan_out[11] : edt_bypass_in[12];
   assign edt_scan_in[13] = edt_bypass ? edt_scan_out[12] : edt_bypass_in[13];
   assign edt_scan_in[14] = edt_bypass ? edt_scan_out[13] : edt_bypass_in[14];
   assign edt_scan_in[15] = edt_bypass ? edt_scan_out[14] : edt_bypass_in[15];
   assign edt_scan_in[16] = edt_bypass ? edt_scan_out[15] : edt_bypass_in[16];
   assign edt_scan_in[17] = edt_bypass ? edt_scan_out[16] : edt_bypass_in[17];
   assign edt_scan_in[18] = edt_bypass ? edt_scan_out[17] : edt_bypass_in[18];
   assign edt_scan_in[19] = edt_bypass ? edt_scan_out[18] : edt_bypass_in[19];
   assign edt_scan_in[20] = edt_bypass ? edt_scan_out[19] : edt_bypass_in[20];
   assign edt_scan_in[21] = edt_bypass ? edt_scan_out[20] : edt_bypass_in[21];
   assign edt_scan_in[22] = edt_bypass ? edt_scan_out[21] : edt_bypass_in[22];
   assign edt_scan_in[23] = edt_bypass ? edt_scan_out[22] : edt_bypass_in[23];
   assign edt_scan_in[24] = edt_bypass ? edt_scan_out[23] : edt_bypass_in[24];
   assign edt_scan_in[25] = edt_bypass ? edt_scan_out[24] : edt_bypass_in[25];
   assign edt_scan_in[26] = edt_bypass ? edt_scan_out[25] : edt_bypass_in[26];
   assign edt_scan_in[27] = edt_bypass ? edt_scan_out[26] : edt_bypass_in[27];
   assign edt_scan_in[28] = edt_bypass ? edt_scan_out[27] : edt_bypass_in[28];
   assign edt_scan_in[29] = edt_bypass ? edt_scan_out[28] : edt_bypass_in[29];
   assign edt_scan_in[30] = edt_bypass ? edt_scan_out[29] : edt_bypass_in[30];
   assign edt_scan_in[31] = edt_bypass ? edt_scan_out[30] : edt_bypass_in[31];
   assign edt_scan_in[32] = edt_bypass ? edt_scan_out[31] : edt_bypass_in[32];
   assign edt_scan_in[33] = edt_bypass ? edt_scan_out[32] : edt_bypass_in[33];
   assign edt_scan_in[34] = edt_bypass ? edt_scan_out[33] : edt_bypass_in[34];
   assign edt_scan_in[35] = edt_bypass ? edt_scan_out[34] : edt_bypass_in[35];
   assign edt_scan_in[36] = edt_bypass ? edt_scan_out[35] : edt_bypass_in[36];
   assign edt_scan_in[37] = edt_bypass ? edt_scan_out[36] : edt_bypass_in[37];
   assign edt_scan_in[38] = edt_bypass ? edt_scan_out[37] : edt_bypass_in[38];
   assign edt_scan_in[39] = edt_bypass ? edt_scan_out[38] : edt_bypass_in[39];
   assign edt_scan_in[40] = edt_bypass ? edt_scan_out[39] : edt_bypass_in[40];
   assign edt_scan_in[41] = edt_bypass ? edt_scan_out[40] : edt_bypass_in[41];
   assign edt_scan_in[42] = edt_bypass ? edt_scan_out[41] : edt_bypass_in[42];
   assign edt_scan_in[43] = edt_bypass ? edt_scan_out[42] : edt_bypass_in[43];
   assign edt_scan_in[44] = edt_bypass ? edt_scan_out[43] : edt_bypass_in[44];
   assign edt_scan_in[45] = edt_bypass ? edt_scan_out[44] : edt_bypass_in[45];
   assign edt_scan_in[46] = edt_bypass ? edt_scan_out[45] : edt_bypass_in[46];
   assign edt_scan_in[47] = edt_bypass ? edt_scan_out[46] : edt_bypass_in[47];
   assign edt_scan_in[48] = edt_bypass ? edt_scan_out[47] : edt_bypass_in[48];
   assign edt_scan_in[49] = edt_bypass ? edt_scan_out[48] : edt_bypass_in[49];
   assign edt_scan_in[50] = edt_bypass ? edt_scan_out[49] : edt_bypass_in[50];
   assign edt_scan_in[51] = edt_bypass ? edt_scan_out[50] : edt_bypass_in[51];
   assign edt_scan_in[52] = edt_bypass ? edt_scan_out[51] : edt_bypass_in[52];
   assign edt_scan_in[53] = edt_bypass ? edt_scan_out[52] : edt_bypass_in[53];
   assign edt_scan_in[54] = edt_bypass ? edt_scan_out[53] : edt_bypass_in[54];
   assign edt_scan_in[55] = edt_bypass ? edt_scan_out[54] : edt_bypass_in[55];
   assign edt_scan_in[56] = edt_bypass ? edt_scan_out[55] : edt_bypass_in[56];
   assign edt_scan_in[57] = edt_bypass ? edt_scan_out[56] : edt_bypass_in[57];
   assign edt_scan_in[58] = edt_bypass ? edt_scan_out[57] : edt_bypass_in[58];
   assign edt_scan_in[59] = edt_bypass ? edt_scan_out[58] : edt_bypass_in[59];
   assign edt_scan_in[60] = edt_bypass ? edt_scan_out[59] : edt_bypass_in[60];
   assign edt_scan_in[61] = edt_bypass ? edt_scan_out[60] : edt_bypass_in[61];
   assign edt_scan_in[62] = edt_bypass ? edt_scan_out[61] : edt_bypass_in[62];
   assign edt_scan_in[63] = edt_bypass ? edt_scan_out[62] : edt_bypass_in[63];
   assign edt_scan_in[64] = edt_bypass ? edt_scan_out[63] : edt_bypass_in[64];
   assign edt_scan_in[65] = edt_bypass ? edt_scan_out[64] : edt_bypass_in[65];
   assign edt_scan_in[66] = edt_bypass ? edt_scan_out[65] : edt_bypass_in[66];
   assign edt_scan_in[67] = edt_bypass ? edt_scan_out[66] : edt_bypass_in[67];
   assign edt_scan_in[68] = edt_bypass ? edt_scan_out[67] : edt_bypass_in[68];
   assign edt_scan_in[69] = edt_bypass ? edt_scan_out[68] : edt_bypass_in[69];
   assign edt_scan_in[70] = edt_bypass ? edt_scan_out[69] : edt_bypass_in[70];
   assign edt_scan_in[71] = edt_bypass ? edt_scan_out[70] : edt_bypass_in[71];
   assign edt_scan_in[72] = edt_bypass ? edt_scan_out[71] : edt_bypass_in[72];
   assign edt_scan_in[73] = edt_bypass ? edt_scan_out[72] : edt_bypass_in[73];
   assign edt_scan_in[74] = edt_bypass ? edt_scan_out[73] : edt_bypass_in[74];
   assign edt_scan_in[75] = edt_bypass ? edt_scan_out[74] : edt_bypass_in[75];
   assign edt_scan_in[76] = edt_bypass ? edt_scan_out[75] : edt_bypass_in[76];
   assign edt_scan_in[77] = edt_bypass ? edt_scan_out[76] : edt_bypass_in[77];
   assign edt_scan_in[78] = edt_bypass ? edt_scan_out[77] : edt_bypass_in[78];
   assign edt_scan_in[79] = edt_bypass ? edt_scan_out[78] : edt_bypass_in[79];
   assign edt_scan_in[80] = edt_bypass ? edt_scan_out[79] : edt_bypass_in[80];
   assign edt_scan_in[81] = edt_bypass ? edt_scan_out[80] : edt_bypass_in[81];
   assign edt_scan_in[82] = edt_bypass ? edt_scan_out[81] : edt_bypass_in[82];
   assign edt_scan_in[83] = edt_bypass ? edt_scan_out[82] : edt_bypass_in[83];
   assign edt_scan_in[84] = edt_bypass ? edt_scan_out[83] : edt_bypass_in[84];
   assign edt_scan_in[85] = edt_bypass ? edt_scan_out[84] : edt_bypass_in[85];
   assign edt_scan_in[86] = edt_bypass ? edt_scan_out[85] : edt_bypass_in[86];
   assign edt_scan_in[87] = edt_bypass ? edt_scan_out[86] : edt_bypass_in[87];
   assign edt_scan_in[88] = edt_bypass ? edt_scan_out[87] : edt_bypass_in[88];
   assign edt_scan_in[89] = edt_bypass ? edt_scan_out[88] : edt_bypass_in[89];
   assign edt_scan_in[90] = edt_bypass ? edt_scan_out[89] : edt_bypass_in[90];
   assign edt_scan_in[91] = edt_bypass ? edt_scan_out[90] : edt_bypass_in[91];
   assign edt_scan_in[92] = edt_bypass ? edt_scan_out[91] : edt_bypass_in[92];
   assign edt_scan_in[93] = edt_bypass ? edt_scan_out[92] : edt_bypass_in[93];
   assign edt_scan_in[94] = edt_bypass ? edt_scan_out[93] : edt_bypass_in[94];
   assign edt_scan_in[95] = edt_bypass ? edt_scan_out[94] : edt_bypass_in[95];
   assign edt_scan_in[96] = edt_bypass ? edt_scan_out[95] : edt_bypass_in[96];
   assign edt_scan_in[97] = edt_bypass ? edt_scan_out[96] : edt_bypass_in[97];
   assign edt_scan_in[98] = edt_bypass ? edt_scan_out[97] : edt_bypass_in[98];
   assign edt_scan_in[99] = edt_bypass ? edt_scan_out[98] : edt_bypass_in[99];
   assign edt_scan_in[100] = edt_bypass ? edt_scan_out[99] : edt_bypass_in[100];
   assign edt_scan_in[101] = edt_bypass ? edt_scan_out[100] : edt_bypass_in[101];
   assign edt_scan_in[102] = edt_bypass ? edt_scan_out[101] : edt_bypass_in[102];
   assign edt_scan_in[103] = edt_bypass ? edt_scan_out[102] : edt_bypass_in[103];
   assign edt_scan_in[104] = edt_bypass ? edt_scan_out[103] : edt_bypass_in[104];
   assign edt_scan_in[105] = edt_bypass ? edt_scan_out[104] : edt_bypass_in[105];
   assign edt_scan_in[106] = edt_bypass ? edt_scan_out[105] : edt_bypass_in[106];
   assign edt_scan_in[107] = edt_bypass ? edt_scan_out[106] : edt_bypass_in[107];
   assign edt_scan_in[108] = edt_bypass ? edt_scan_out[107] : edt_bypass_in[108];
   assign edt_scan_in[109] = edt_bypass ? edt_scan_out[108] : edt_bypass_in[109];
   assign edt_scan_in[110] = edt_bypass ? edt_scan_out[109] : edt_bypass_in[110];
   assign edt_scan_in[111] = edt_bypass ? edt_scan_out[110] : edt_bypass_in[111];
   assign edt_scan_in[112] = edt_bypass ? edt_scan_out[111] : edt_bypass_in[112];
   assign edt_scan_in[113] = edt_bypass ? edt_scan_out[112] : edt_bypass_in[113];
   assign edt_scan_in[114] = edt_bypass ? edt_scan_out[113] : edt_bypass_in[114];
   assign edt_scan_in[115] = edt_bypass ? edt_scan_out[114] : edt_bypass_in[115];
   assign edt_scan_in[116] = edt_bypass ? edt_scan_out[115] : edt_bypass_in[116];
   assign edt_scan_in[117] = edt_bypass ? edt_scan_out[116] : edt_bypass_in[117];
   assign edt_scan_in[118] = edt_bypass ? edt_scan_out[117] : edt_bypass_in[118];
   assign edt_scan_in[119] = edt_bypass ? edt_scan_out[118] : edt_bypass_in[119];
   assign edt_scan_in[120] = edt_bypass ? edt_scan_out[119] : edt_bypass_in[120];
   assign edt_scan_in[121] = edt_bypass ? edt_scan_out[120] : edt_bypass_in[121];
   assign edt_scan_in[122] = edt_bypass ? edt_scan_out[121] : edt_bypass_in[122];
   assign edt_scan_in[123] = edt_bypass ? edt_scan_out[122] : edt_bypass_in[123];
   assign edt_scan_in[124] = edt_bypass ? edt_scan_out[123] : edt_bypass_in[124];
   assign edt_scan_in[125] = edt_bypass ? edt_scan_out[124] : edt_bypass_in[125];
   assign edt_scan_in[126] = edt_bypass ? edt_scan_out[125] : edt_bypass_in[126];
   assign edt_scan_in[127] = edt_bypass ? edt_scan_out[126] : edt_bypass_in[127];
   assign edt_scan_in[128] = edt_bypass ? edt_scan_out[127] : edt_bypass_in[128];
   assign edt_scan_in[129] = edt_bypass ? edt_scan_out[128] : edt_bypass_in[129];
   assign edt_scan_in[130] = edt_bypass ? edt_scan_out[129] : edt_bypass_in[130];
   assign edt_scan_in[131] = edt_bypass ? edt_scan_out[130] : edt_bypass_in[131];
   assign edt_scan_in[132] = edt_bypass ? edt_scan_out[131] : edt_bypass_in[132];
   assign edt_scan_in[133] = edt_bypass ? edt_scan_out[132] : edt_bypass_in[133];
   assign edt_scan_in[134] = edt_bypass ? edt_scan_out[133] : edt_bypass_in[134];
   assign edt_scan_in[135] = edt_bypass ? edt_scan_out[134] : edt_bypass_in[135];
   assign edt_scan_in[136] = edt_bypass ? edt_scan_out[135] : edt_bypass_in[136];
   assign edt_scan_in[137] = edt_bypass ? edt_scan_out[136] : edt_bypass_in[137];
   assign edt_scan_in[138] = edt_bypass ? edt_scan_out[137] : edt_bypass_in[138];
   assign edt_scan_in[139] = edt_bypass ? edt_scan_out[138] : edt_bypass_in[139];
   assign edt_scan_in[140] = edt_bypass ? edt_scan_out[139] : edt_bypass_in[140];
   assign edt_scan_in[141] = edt_bypass ? edt_scan_out[140] : edt_bypass_in[141];
   assign edt_scan_in[142] = edt_bypass ? edt_scan_out[141] : edt_bypass_in[142];
   assign edt_scan_in[143] = edt_bypass ? edt_scan_out[142] : edt_bypass_in[143];
   assign edt_scan_in[144] = edt_bypass ? edt_scan_out[143] : edt_bypass_in[144];
   assign edt_scan_in[145] = edt_bypass ? edt_scan_out[144] : edt_bypass_in[145];
   assign edt_scan_in[146] = edt_bypass ? edt_scan_out[145] : edt_bypass_in[146];
   assign edt_scan_in[147] = edt_bypass ? edt_scan_out[146] : edt_bypass_in[147];
   assign edt_scan_in[148] = edt_bypass ? edt_scan_out[147] : edt_bypass_in[148];
   assign edt_scan_in[149] = edt_bypass ? edt_scan_out[148] : edt_bypass_in[149];
   assign edt_scan_in[150] = edt_bypass ? edt_scan_out[149] : edt_bypass_in[150];
   assign edt_scan_in[151] = edt_bypass ? edt_scan_out[150] : edt_bypass_in[151];
   assign edt_scan_in[152] = edt_bypass ? edt_scan_out[151] : edt_bypass_in[152];
   assign edt_scan_in[153] = edt_bypass ? edt_scan_out[152] : edt_bypass_in[153];
   assign edt_scan_in[154] = edt_bypass ? edt_scan_out[153] : edt_bypass_in[154];
   assign edt_scan_in[155] = edt_bypass ? edt_scan_out[154] : edt_bypass_in[155];
   assign edt_scan_in[156] = edt_bypass ? edt_scan_out[155] : edt_bypass_in[156];
   assign edt_scan_in[157] = edt_bypass ? edt_scan_out[156] : edt_bypass_in[157];
   assign edt_scan_in[158] = edt_bypass ? edt_scan_out[157] : edt_bypass_in[158];
   assign edt_scan_in[159] = edt_bypass ? edt_scan_out[158] : edt_bypass_in[159];
   assign edt_scan_in[160] = edt_bypass ? edt_scan_out[159] : edt_bypass_in[160];
   assign edt_scan_in[161] = edt_bypass ? edt_scan_out[160] : edt_bypass_in[161];
   assign edt_scan_in[162] = edt_bypass ? edt_scan_out[161] : edt_bypass_in[162];
   assign edt_scan_in[163] = edt_bypass ? edt_scan_out[162] : edt_bypass_in[163];
   assign edt_scan_in[164] = edt_bypass ? edt_scan_out[163] : edt_bypass_in[164];
   assign edt_scan_in[165] = edt_bypass ? edt_scan_out[164] : edt_bypass_in[165];
   assign edt_scan_in[166] = edt_bypass ? edt_scan_out[165] : edt_bypass_in[166];
   assign edt_scan_in[167] = edt_bypass ? edt_scan_out[166] : edt_bypass_in[167];
   assign edt_scan_in[168] = edt_bypass ? edt_scan_out[167] : edt_bypass_in[168];
   assign edt_scan_in[169] = edt_bypass ? edt_scan_out[168] : edt_bypass_in[169];
   assign edt_scan_in[170] = edt_bypass ? edt_scan_out[169] : edt_bypass_in[170];
   assign edt_scan_in[171] = edt_bypass ? edt_scan_out[170] : edt_bypass_in[171];
   assign edt_scan_in[172] = edt_bypass ? edt_scan_out[171] : edt_bypass_in[172];
   assign edt_scan_in[173] = edt_bypass ? edt_scan_out[172] : edt_bypass_in[173];
   assign edt_scan_in[174] = edt_bypass ? edt_scan_out[173] : edt_bypass_in[174];
   assign edt_scan_in[175] = edt_bypass ? edt_scan_out[174] : edt_bypass_in[175];
   assign edt_scan_in[176] = edt_bypass ? edt_scan_out[175] : edt_bypass_in[176];
   assign edt_scan_in[177] = edt_bypass ? edt_scan_out[176] : edt_bypass_in[177];
   assign edt_scan_in[178] = edt_bypass ? edt_scan_out[177] : edt_bypass_in[178];
   assign edt_scan_in[179] = edt_bypass ? edt_scan_out[178] : edt_bypass_in[179];
   assign edt_scan_in[180] = edt_bypass ? edt_scan_out[179] : edt_bypass_in[180];
   assign edt_scan_in[181] = edt_bypass ? edt_scan_out[180] : edt_bypass_in[181];
   assign edt_scan_in[182] = edt_bypass ? edt_scan_out[181] : edt_bypass_in[182];
   assign edt_scan_in[183] = edt_bypass ? edt_scan_out[182] : edt_bypass_in[183];
   assign edt_scan_in[184] = edt_bypass ? edt_scan_out[183] : edt_bypass_in[184];
   assign edt_scan_in[185] = edt_bypass ? edt_scan_out[184] : edt_bypass_in[185];
   assign edt_scan_in[186] = edt_bypass ? edt_channels_in[1] : edt_bypass_in[186];
   assign edt_scan_in[187] = edt_bypass ? edt_scan_out[186] : edt_bypass_in[187];
   assign edt_scan_in[188] = edt_bypass ? edt_scan_out[187] : edt_bypass_in[188];
   assign edt_scan_in[189] = edt_bypass ? edt_scan_out[188] : edt_bypass_in[189];
   assign edt_scan_in[190] = edt_bypass ? edt_scan_out[189] : edt_bypass_in[190];
   assign edt_scan_in[191] = edt_bypass ? edt_scan_out[190] : edt_bypass_in[191];
   assign edt_scan_in[192] = edt_bypass ? edt_scan_out[191] : edt_bypass_in[192];
   assign edt_scan_in[193] = edt_bypass ? edt_scan_out[192] : edt_bypass_in[193];
   assign edt_scan_in[194] = edt_bypass ? edt_scan_out[193] : edt_bypass_in[194];
   assign edt_scan_in[195] = edt_bypass ? edt_scan_out[194] : edt_bypass_in[195];
   assign edt_scan_in[196] = edt_bypass ? edt_scan_out[195] : edt_bypass_in[196];
   assign edt_scan_in[197] = edt_bypass ? edt_scan_out[196] : edt_bypass_in[197];
   assign edt_scan_in[198] = edt_bypass ? edt_scan_out[197] : edt_bypass_in[198];
   assign edt_scan_in[199] = edt_bypass ? edt_scan_out[198] : edt_bypass_in[199];
   assign edt_scan_in[200] = edt_bypass ? edt_scan_out[199] : edt_bypass_in[200];
   assign edt_scan_in[201] = edt_bypass ? edt_scan_out[200] : edt_bypass_in[201];
   assign edt_scan_in[202] = edt_bypass ? edt_scan_out[201] : edt_bypass_in[202];
   assign edt_scan_in[203] = edt_bypass ? edt_scan_out[202] : edt_bypass_in[203];
   assign edt_scan_in[204] = edt_bypass ? edt_scan_out[203] : edt_bypass_in[204];
   assign edt_scan_in[205] = edt_bypass ? edt_scan_out[204] : edt_bypass_in[205];
   assign edt_scan_in[206] = edt_bypass ? edt_scan_out[205] : edt_bypass_in[206];
   assign edt_scan_in[207] = edt_bypass ? edt_scan_out[206] : edt_bypass_in[207];
   assign edt_scan_in[208] = edt_bypass ? edt_scan_out[207] : edt_bypass_in[208];
   assign edt_scan_in[209] = edt_bypass ? edt_scan_out[208] : edt_bypass_in[209];
   assign edt_scan_in[210] = edt_bypass ? edt_scan_out[209] : edt_bypass_in[210];
   assign edt_scan_in[211] = edt_bypass ? edt_scan_out[210] : edt_bypass_in[211];
   assign edt_scan_in[212] = edt_bypass ? edt_scan_out[211] : edt_bypass_in[212];
   assign edt_scan_in[213] = edt_bypass ? edt_scan_out[212] : edt_bypass_in[213];
   assign edt_scan_in[214] = edt_bypass ? edt_scan_out[213] : edt_bypass_in[214];
   assign edt_scan_in[215] = edt_bypass ? edt_scan_out[214] : edt_bypass_in[215];
   assign edt_scan_in[216] = edt_bypass ? edt_scan_out[215] : edt_bypass_in[216];
   assign edt_scan_in[217] = edt_bypass ? edt_scan_out[216] : edt_bypass_in[217];
   assign edt_scan_in[218] = edt_bypass ? edt_scan_out[217] : edt_bypass_in[218];
   assign edt_scan_in[219] = edt_bypass ? edt_scan_out[218] : edt_bypass_in[219];
   assign edt_scan_in[220] = edt_bypass ? edt_scan_out[219] : edt_bypass_in[220];
   assign edt_scan_in[221] = edt_bypass ? edt_scan_out[220] : edt_bypass_in[221];
   assign edt_scan_in[222] = edt_bypass ? edt_scan_out[221] : edt_bypass_in[222];
   assign edt_scan_in[223] = edt_bypass ? edt_scan_out[222] : edt_bypass_in[223];
   assign edt_scan_in[224] = edt_bypass ? edt_scan_out[223] : edt_bypass_in[224];
   assign edt_scan_in[225] = edt_bypass ? edt_scan_out[224] : edt_bypass_in[225];
   assign edt_scan_in[226] = edt_bypass ? edt_scan_out[225] : edt_bypass_in[226];
   assign edt_scan_in[227] = edt_bypass ? edt_scan_out[226] : edt_bypass_in[227];
   assign edt_scan_in[228] = edt_bypass ? edt_scan_out[227] : edt_bypass_in[228];
   assign edt_scan_in[229] = edt_bypass ? edt_scan_out[228] : edt_bypass_in[229];
   assign edt_scan_in[230] = edt_bypass ? edt_scan_out[229] : edt_bypass_in[230];
   assign edt_scan_in[231] = edt_bypass ? edt_scan_out[230] : edt_bypass_in[231];
   assign edt_scan_in[232] = edt_bypass ? edt_scan_out[231] : edt_bypass_in[232];
   assign edt_scan_in[233] = edt_bypass ? edt_scan_out[232] : edt_bypass_in[233];
   assign edt_scan_in[234] = edt_bypass ? edt_scan_out[233] : edt_bypass_in[234];
   assign edt_scan_in[235] = edt_bypass ? edt_scan_out[234] : edt_bypass_in[235];
   assign edt_scan_in[236] = edt_bypass ? edt_scan_out[235] : edt_bypass_in[236];
   assign edt_scan_in[237] = edt_bypass ? edt_scan_out[236] : edt_bypass_in[237];
   assign edt_scan_in[238] = edt_bypass ? edt_scan_out[237] : edt_bypass_in[238];
   assign edt_scan_in[239] = edt_bypass ? edt_scan_out[238] : edt_bypass_in[239];
   assign edt_scan_in[240] = edt_bypass ? edt_scan_out[239] : edt_bypass_in[240];
   assign edt_scan_in[241] = edt_bypass ? edt_scan_out[240] : edt_bypass_in[241];
   assign edt_scan_in[242] = edt_bypass ? edt_scan_out[241] : edt_bypass_in[242];
   assign edt_scan_in[243] = edt_bypass ? edt_scan_out[242] : edt_bypass_in[243];
   assign edt_scan_in[244] = edt_bypass ? edt_scan_out[243] : edt_bypass_in[244];
   assign edt_scan_in[245] = edt_bypass ? edt_scan_out[244] : edt_bypass_in[245];
   assign edt_scan_in[246] = edt_bypass ? edt_scan_out[245] : edt_bypass_in[246];
   assign edt_scan_in[247] = edt_bypass ? edt_scan_out[246] : edt_bypass_in[247];
   assign edt_scan_in[248] = edt_bypass ? edt_scan_out[247] : edt_bypass_in[248];
   assign edt_scan_in[249] = edt_bypass ? edt_scan_out[248] : edt_bypass_in[249];
   assign edt_scan_in[250] = edt_bypass ? edt_scan_out[249] : edt_bypass_in[250];
   assign edt_scan_in[251] = edt_bypass ? edt_scan_out[250] : edt_bypass_in[251];
   assign edt_scan_in[252] = edt_bypass ? edt_scan_out[251] : edt_bypass_in[252];
   assign edt_scan_in[253] = edt_bypass ? edt_scan_out[252] : edt_bypass_in[253];
   assign edt_scan_in[254] = edt_bypass ? edt_scan_out[253] : edt_bypass_in[254];
   assign edt_scan_in[255] = edt_bypass ? edt_scan_out[254] : edt_bypass_in[255];
   assign edt_scan_in[256] = edt_bypass ? edt_scan_out[255] : edt_bypass_in[256];
   assign edt_scan_in[257] = edt_bypass ? edt_scan_out[256] : edt_bypass_in[257];
   assign edt_scan_in[258] = edt_bypass ? edt_scan_out[257] : edt_bypass_in[258];
   assign edt_scan_in[259] = edt_bypass ? edt_scan_out[258] : edt_bypass_in[259];
   assign edt_scan_in[260] = edt_bypass ? edt_scan_out[259] : edt_bypass_in[260];
   assign edt_scan_in[261] = edt_bypass ? edt_scan_out[260] : edt_bypass_in[261];
   assign edt_scan_in[262] = edt_bypass ? edt_scan_out[261] : edt_bypass_in[262];
   assign edt_scan_in[263] = edt_bypass ? edt_scan_out[262] : edt_bypass_in[263];
   assign edt_scan_in[264] = edt_bypass ? edt_scan_out[263] : edt_bypass_in[264];
   assign edt_scan_in[265] = edt_bypass ? edt_scan_out[264] : edt_bypass_in[265];
   assign edt_scan_in[266] = edt_bypass ? edt_scan_out[265] : edt_bypass_in[266];
   assign edt_scan_in[267] = edt_bypass ? edt_scan_out[266] : edt_bypass_in[267];
   assign edt_scan_in[268] = edt_bypass ? edt_scan_out[267] : edt_bypass_in[268];
   assign edt_scan_in[269] = edt_bypass ? edt_scan_out[268] : edt_bypass_in[269];
   assign edt_scan_in[270] = edt_bypass ? edt_scan_out[269] : edt_bypass_in[270];
   assign edt_scan_in[271] = edt_bypass ? edt_scan_out[270] : edt_bypass_in[271];
   assign edt_scan_in[272] = edt_bypass ? edt_scan_out[271] : edt_bypass_in[272];
   assign edt_scan_in[273] = edt_bypass ? edt_scan_out[272] : edt_bypass_in[273];
   assign edt_scan_in[274] = edt_bypass ? edt_scan_out[273] : edt_bypass_in[274];
   assign edt_scan_in[275] = edt_bypass ? edt_scan_out[274] : edt_bypass_in[275];
   assign edt_scan_in[276] = edt_bypass ? edt_scan_out[275] : edt_bypass_in[276];
   assign edt_scan_in[277] = edt_bypass ? edt_scan_out[276] : edt_bypass_in[277];
   assign edt_scan_in[278] = edt_bypass ? edt_scan_out[277] : edt_bypass_in[278];
   assign edt_scan_in[279] = edt_bypass ? edt_scan_out[278] : edt_bypass_in[279];
   assign edt_scan_in[280] = edt_bypass ? edt_scan_out[279] : edt_bypass_in[280];
   assign edt_scan_in[281] = edt_bypass ? edt_scan_out[280] : edt_bypass_in[281];
   assign edt_scan_in[282] = edt_bypass ? edt_scan_out[281] : edt_bypass_in[282];
   assign edt_scan_in[283] = edt_bypass ? edt_scan_out[282] : edt_bypass_in[283];
   assign edt_scan_in[284] = edt_bypass ? edt_scan_out[283] : edt_bypass_in[284];
   assign edt_scan_in[285] = edt_bypass ? edt_scan_out[284] : edt_bypass_in[285];
   assign edt_scan_in[286] = edt_bypass ? edt_scan_out[285] : edt_bypass_in[286];
   assign edt_scan_in[287] = edt_bypass ? edt_scan_out[286] : edt_bypass_in[287];
   assign edt_scan_in[288] = edt_bypass ? edt_scan_out[287] : edt_bypass_in[288];
   assign edt_scan_in[289] = edt_bypass ? edt_scan_out[288] : edt_bypass_in[289];
   assign edt_scan_in[290] = edt_bypass ? edt_scan_out[289] : edt_bypass_in[290];
   assign edt_scan_in[291] = edt_bypass ? edt_scan_out[290] : edt_bypass_in[291];
   assign edt_scan_in[292] = edt_bypass ? edt_scan_out[291] : edt_bypass_in[292];
   assign edt_scan_in[293] = edt_bypass ? edt_scan_out[292] : edt_bypass_in[293];
   assign edt_scan_in[294] = edt_bypass ? edt_scan_out[293] : edt_bypass_in[294];
   assign edt_scan_in[295] = edt_bypass ? edt_scan_out[294] : edt_bypass_in[295];
   assign edt_scan_in[296] = edt_bypass ? edt_scan_out[295] : edt_bypass_in[296];
   assign edt_scan_in[297] = edt_bypass ? edt_scan_out[296] : edt_bypass_in[297];
   assign edt_scan_in[298] = edt_bypass ? edt_scan_out[297] : edt_bypass_in[298];
   assign edt_scan_in[299] = edt_bypass ? edt_scan_out[298] : edt_bypass_in[299];
   assign edt_scan_in[300] = edt_bypass ? edt_scan_out[299] : edt_bypass_in[300];
   assign edt_scan_in[301] = edt_bypass ? edt_scan_out[300] : edt_bypass_in[301];
   assign edt_scan_in[302] = edt_bypass ? edt_scan_out[301] : edt_bypass_in[302];
   assign edt_scan_in[303] = edt_bypass ? edt_scan_out[302] : edt_bypass_in[303];
   assign edt_scan_in[304] = edt_bypass ? edt_scan_out[303] : edt_bypass_in[304];
   assign edt_scan_in[305] = edt_bypass ? edt_scan_out[304] : edt_bypass_in[305];
   assign edt_scan_in[306] = edt_bypass ? edt_scan_out[305] : edt_bypass_in[306];
   assign edt_scan_in[307] = edt_bypass ? edt_scan_out[306] : edt_bypass_in[307];
   assign edt_scan_in[308] = edt_bypass ? edt_scan_out[307] : edt_bypass_in[308];
   assign edt_scan_in[309] = edt_bypass ? edt_scan_out[308] : edt_bypass_in[309];
   assign edt_scan_in[310] = edt_bypass ? edt_scan_out[309] : edt_bypass_in[310];
   assign edt_scan_in[311] = edt_bypass ? edt_scan_out[310] : edt_bypass_in[311];
   assign edt_scan_in[312] = edt_bypass ? edt_scan_out[311] : edt_bypass_in[312];
   assign edt_scan_in[313] = edt_bypass ? edt_scan_out[312] : edt_bypass_in[313];
   assign edt_scan_in[314] = edt_bypass ? edt_scan_out[313] : edt_bypass_in[314];
   assign edt_scan_in[315] = edt_bypass ? edt_scan_out[314] : edt_bypass_in[315];
   assign edt_scan_in[316] = edt_bypass ? edt_scan_out[315] : edt_bypass_in[316];
   assign edt_scan_in[317] = edt_bypass ? edt_scan_out[316] : edt_bypass_in[317];
   assign edt_scan_in[318] = edt_bypass ? edt_scan_out[317] : edt_bypass_in[318];
   assign edt_scan_in[319] = edt_bypass ? edt_scan_out[318] : edt_bypass_in[319];
   assign edt_scan_in[320] = edt_bypass ? edt_scan_out[319] : edt_bypass_in[320];
   assign edt_scan_in[321] = edt_bypass ? edt_scan_out[320] : edt_bypass_in[321];
   assign edt_scan_in[322] = edt_bypass ? edt_scan_out[321] : edt_bypass_in[322];
   assign edt_scan_in[323] = edt_bypass ? edt_scan_out[322] : edt_bypass_in[323];
   assign edt_scan_in[324] = edt_bypass ? edt_scan_out[323] : edt_bypass_in[324];
   assign edt_scan_in[325] = edt_bypass ? edt_scan_out[324] : edt_bypass_in[325];
   assign edt_scan_in[326] = edt_bypass ? edt_scan_out[325] : edt_bypass_in[326];
   assign edt_scan_in[327] = edt_bypass ? edt_scan_out[326] : edt_bypass_in[327];
   assign edt_scan_in[328] = edt_bypass ? edt_scan_out[327] : edt_bypass_in[328];
   assign edt_scan_in[329] = edt_bypass ? edt_scan_out[328] : edt_bypass_in[329];
   assign edt_scan_in[330] = edt_bypass ? edt_scan_out[329] : edt_bypass_in[330];
   assign edt_scan_in[331] = edt_bypass ? edt_scan_out[330] : edt_bypass_in[331];
   assign edt_scan_in[332] = edt_bypass ? edt_scan_out[331] : edt_bypass_in[332];
   assign edt_scan_in[333] = edt_bypass ? edt_scan_out[332] : edt_bypass_in[333];
   assign edt_scan_in[334] = edt_bypass ? edt_scan_out[333] : edt_bypass_in[334];
   assign edt_scan_in[335] = edt_bypass ? edt_scan_out[334] : edt_bypass_in[335];
   assign edt_scan_in[336] = edt_bypass ? edt_scan_out[335] : edt_bypass_in[336];
   assign edt_scan_in[337] = edt_bypass ? edt_scan_out[336] : edt_bypass_in[337];
   assign edt_scan_in[338] = edt_bypass ? edt_scan_out[337] : edt_bypass_in[338];
   assign edt_scan_in[339] = edt_bypass ? edt_scan_out[338] : edt_bypass_in[339];
   assign edt_scan_in[340] = edt_bypass ? edt_scan_out[339] : edt_bypass_in[340];
   assign edt_scan_in[341] = edt_bypass ? edt_scan_out[340] : edt_bypass_in[341];
   assign edt_scan_in[342] = edt_bypass ? edt_scan_out[341] : edt_bypass_in[342];
   assign edt_scan_in[343] = edt_bypass ? edt_scan_out[342] : edt_bypass_in[343];
   assign edt_scan_in[344] = edt_bypass ? edt_scan_out[343] : edt_bypass_in[344];
   assign edt_scan_in[345] = edt_bypass ? edt_scan_out[344] : edt_bypass_in[345];
   assign edt_scan_in[346] = edt_bypass ? edt_scan_out[345] : edt_bypass_in[346];
   assign edt_scan_in[347] = edt_bypass ? edt_scan_out[346] : edt_bypass_in[347];
   assign edt_scan_in[348] = edt_bypass ? edt_scan_out[347] : edt_bypass_in[348];
   assign edt_scan_in[349] = edt_bypass ? edt_scan_out[348] : edt_bypass_in[349];
   assign edt_scan_in[350] = edt_bypass ? edt_scan_out[349] : edt_bypass_in[350];
   assign edt_scan_in[351] = edt_bypass ? edt_scan_out[350] : edt_bypass_in[351];
   assign edt_scan_in[352] = edt_bypass ? edt_scan_out[351] : edt_bypass_in[352];
   assign edt_scan_in[353] = edt_bypass ? edt_scan_out[352] : edt_bypass_in[353];
   assign edt_scan_in[354] = edt_bypass ? edt_scan_out[353] : edt_bypass_in[354];
   assign edt_scan_in[355] = edt_bypass ? edt_scan_out[354] : edt_bypass_in[355];
   assign edt_scan_in[356] = edt_bypass ? edt_scan_out[355] : edt_bypass_in[356];
   assign edt_scan_in[357] = edt_bypass ? edt_scan_out[356] : edt_bypass_in[357];
   assign edt_scan_in[358] = edt_bypass ? edt_scan_out[357] : edt_bypass_in[358];
   assign edt_scan_in[359] = edt_bypass ? edt_scan_out[358] : edt_bypass_in[359];
   assign edt_scan_in[360] = edt_bypass ? edt_scan_out[359] : edt_bypass_in[360];
   assign edt_scan_in[361] = edt_bypass ? edt_scan_out[360] : edt_bypass_in[361];
   assign edt_scan_in[362] = edt_bypass ? edt_scan_out[361] : edt_bypass_in[362];
   assign edt_scan_in[363] = edt_bypass ? edt_scan_out[362] : edt_bypass_in[363];
   assign edt_scan_in[364] = edt_bypass ? edt_scan_out[363] : edt_bypass_in[364];
   assign edt_scan_in[365] = edt_bypass ? edt_scan_out[364] : edt_bypass_in[365];
   assign edt_scan_in[366] = edt_bypass ? edt_scan_out[365] : edt_bypass_in[366];
   assign edt_scan_in[367] = edt_bypass ? edt_scan_out[366] : edt_bypass_in[367];
   assign edt_scan_in[368] = edt_bypass ? edt_scan_out[367] : edt_bypass_in[368];
   assign edt_scan_in[369] = edt_bypass ? edt_scan_out[368] : edt_bypass_in[369];
   assign edt_scan_in[370] = edt_bypass ? edt_scan_out[369] : edt_bypass_in[370];

   assign edt_channels_out[0] = edt_bypass ? edt_scan_out[185] : edt_bypass_out[0];
   assign edt_channels_out[1] = edt_bypass ? edt_scan_out[370] : edt_bypass_out[1];
endmodule


module firebird7_in_gate2_tessent_edt_intest_edt (
   input  wire         edt_clock,
   input  wire         edt_update,
   input  wire         edt_low_power_shift_en,
   input  wire         edt_bypass,
   input  wire [  3:0] edt_channels_in,
   output wire [  1:0] edt_channels_out,
   output wire [370:0] edt_scan_in,
   input  wire [370:0] edt_scan_out
);
   wire   [370:0] edt_decompressor_out;
   wire   [370:0] edt_bypass_in;
   wire   [  1:0] edt_bypass_out;
   wire   [185:0] masks_for_compactor_0;
   wire   [184:0] masks_for_compactor_1;
   wire   [  3:0] edt_channels_out_from_controller;
   wire           edt_clock_buf_out;
   wire           edt_update_buf_out;
   wire           edt_bypass_buf_out;
   wire           edt_low_power_shift_en_buf_out;
   wire   [  3:0] edt_channels_in_buf_out;
   wire   [  1:0] edt_channels_out_buf_in;
   wire   [370:0] edt_scan_in_buf_in;
   wire   [370:0] edt_scan_out_buf_out;

   i0scbf000ab1n02x5 tessent_persistent_cell_edt_clock_buf (.clk(edt_clock),
                                                            .clkout(edt_clock_buf_out));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_update_buf (.a(edt_update),
                                                             .o(edt_update_buf_out));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_bypass_buf (.a(edt_bypass),
                                                             .o(edt_bypass_buf_out));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_low_power_shift_en_buf (.a(edt_low_power_shift_en),
                                                                         .o(edt_low_power_shift_en_buf_out));

   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_in_0_buf (.a(edt_channels_in[0]),
                                                                    .o(edt_channels_in_buf_out[0]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_in_1_buf (.a(edt_channels_in[1]),
                                                                    .o(edt_channels_in_buf_out[1]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_in_2_buf (.a(edt_channels_in[2]),
                                                                    .o(edt_channels_in_buf_out[2]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_in_3_buf (.a(edt_channels_in[3]),
                                                                    .o(edt_channels_in_buf_out[3]));

   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_out_0_buf (.a(edt_channels_out_buf_in[0]),
                                                                     .o(edt_channels_out[0]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_channels_out_1_buf (.a(edt_channels_out_buf_in[1]),
                                                                     .o(edt_channels_out[1]));

   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_0_buf (.a(edt_scan_in_buf_in[0]),
                                                                .o(edt_scan_in[0]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_1_buf (.a(edt_scan_in_buf_in[1]),
                                                                .o(edt_scan_in[1]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_2_buf (.a(edt_scan_in_buf_in[2]),
                                                                .o(edt_scan_in[2]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_3_buf (.a(edt_scan_in_buf_in[3]),
                                                                .o(edt_scan_in[3]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_4_buf (.a(edt_scan_in_buf_in[4]),
                                                                .o(edt_scan_in[4]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_5_buf (.a(edt_scan_in_buf_in[5]),
                                                                .o(edt_scan_in[5]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_6_buf (.a(edt_scan_in_buf_in[6]),
                                                                .o(edt_scan_in[6]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_7_buf (.a(edt_scan_in_buf_in[7]),
                                                                .o(edt_scan_in[7]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_8_buf (.a(edt_scan_in_buf_in[8]),
                                                                .o(edt_scan_in[8]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_9_buf (.a(edt_scan_in_buf_in[9]),
                                                                .o(edt_scan_in[9]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_10_buf (.a(edt_scan_in_buf_in[10]),
                                                                 .o(edt_scan_in[10]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_11_buf (.a(edt_scan_in_buf_in[11]),
                                                                 .o(edt_scan_in[11]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_12_buf (.a(edt_scan_in_buf_in[12]),
                                                                 .o(edt_scan_in[12]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_13_buf (.a(edt_scan_in_buf_in[13]),
                                                                 .o(edt_scan_in[13]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_14_buf (.a(edt_scan_in_buf_in[14]),
                                                                 .o(edt_scan_in[14]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_15_buf (.a(edt_scan_in_buf_in[15]),
                                                                 .o(edt_scan_in[15]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_16_buf (.a(edt_scan_in_buf_in[16]),
                                                                 .o(edt_scan_in[16]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_17_buf (.a(edt_scan_in_buf_in[17]),
                                                                 .o(edt_scan_in[17]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_18_buf (.a(edt_scan_in_buf_in[18]),
                                                                 .o(edt_scan_in[18]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_19_buf (.a(edt_scan_in_buf_in[19]),
                                                                 .o(edt_scan_in[19]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_20_buf (.a(edt_scan_in_buf_in[20]),
                                                                 .o(edt_scan_in[20]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_21_buf (.a(edt_scan_in_buf_in[21]),
                                                                 .o(edt_scan_in[21]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_22_buf (.a(edt_scan_in_buf_in[22]),
                                                                 .o(edt_scan_in[22]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_23_buf (.a(edt_scan_in_buf_in[23]),
                                                                 .o(edt_scan_in[23]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_24_buf (.a(edt_scan_in_buf_in[24]),
                                                                 .o(edt_scan_in[24]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_25_buf (.a(edt_scan_in_buf_in[25]),
                                                                 .o(edt_scan_in[25]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_26_buf (.a(edt_scan_in_buf_in[26]),
                                                                 .o(edt_scan_in[26]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_27_buf (.a(edt_scan_in_buf_in[27]),
                                                                 .o(edt_scan_in[27]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_28_buf (.a(edt_scan_in_buf_in[28]),
                                                                 .o(edt_scan_in[28]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_29_buf (.a(edt_scan_in_buf_in[29]),
                                                                 .o(edt_scan_in[29]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_30_buf (.a(edt_scan_in_buf_in[30]),
                                                                 .o(edt_scan_in[30]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_31_buf (.a(edt_scan_in_buf_in[31]),
                                                                 .o(edt_scan_in[31]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_32_buf (.a(edt_scan_in_buf_in[32]),
                                                                 .o(edt_scan_in[32]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_33_buf (.a(edt_scan_in_buf_in[33]),
                                                                 .o(edt_scan_in[33]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_34_buf (.a(edt_scan_in_buf_in[34]),
                                                                 .o(edt_scan_in[34]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_35_buf (.a(edt_scan_in_buf_in[35]),
                                                                 .o(edt_scan_in[35]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_36_buf (.a(edt_scan_in_buf_in[36]),
                                                                 .o(edt_scan_in[36]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_37_buf (.a(edt_scan_in_buf_in[37]),
                                                                 .o(edt_scan_in[37]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_38_buf (.a(edt_scan_in_buf_in[38]),
                                                                 .o(edt_scan_in[38]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_39_buf (.a(edt_scan_in_buf_in[39]),
                                                                 .o(edt_scan_in[39]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_40_buf (.a(edt_scan_in_buf_in[40]),
                                                                 .o(edt_scan_in[40]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_41_buf (.a(edt_scan_in_buf_in[41]),
                                                                 .o(edt_scan_in[41]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_42_buf (.a(edt_scan_in_buf_in[42]),
                                                                 .o(edt_scan_in[42]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_43_buf (.a(edt_scan_in_buf_in[43]),
                                                                 .o(edt_scan_in[43]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_44_buf (.a(edt_scan_in_buf_in[44]),
                                                                 .o(edt_scan_in[44]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_45_buf (.a(edt_scan_in_buf_in[45]),
                                                                 .o(edt_scan_in[45]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_46_buf (.a(edt_scan_in_buf_in[46]),
                                                                 .o(edt_scan_in[46]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_47_buf (.a(edt_scan_in_buf_in[47]),
                                                                 .o(edt_scan_in[47]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_48_buf (.a(edt_scan_in_buf_in[48]),
                                                                 .o(edt_scan_in[48]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_49_buf (.a(edt_scan_in_buf_in[49]),
                                                                 .o(edt_scan_in[49]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_50_buf (.a(edt_scan_in_buf_in[50]),
                                                                 .o(edt_scan_in[50]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_51_buf (.a(edt_scan_in_buf_in[51]),
                                                                 .o(edt_scan_in[51]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_52_buf (.a(edt_scan_in_buf_in[52]),
                                                                 .o(edt_scan_in[52]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_53_buf (.a(edt_scan_in_buf_in[53]),
                                                                 .o(edt_scan_in[53]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_54_buf (.a(edt_scan_in_buf_in[54]),
                                                                 .o(edt_scan_in[54]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_55_buf (.a(edt_scan_in_buf_in[55]),
                                                                 .o(edt_scan_in[55]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_56_buf (.a(edt_scan_in_buf_in[56]),
                                                                 .o(edt_scan_in[56]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_57_buf (.a(edt_scan_in_buf_in[57]),
                                                                 .o(edt_scan_in[57]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_58_buf (.a(edt_scan_in_buf_in[58]),
                                                                 .o(edt_scan_in[58]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_59_buf (.a(edt_scan_in_buf_in[59]),
                                                                 .o(edt_scan_in[59]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_60_buf (.a(edt_scan_in_buf_in[60]),
                                                                 .o(edt_scan_in[60]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_61_buf (.a(edt_scan_in_buf_in[61]),
                                                                 .o(edt_scan_in[61]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_62_buf (.a(edt_scan_in_buf_in[62]),
                                                                 .o(edt_scan_in[62]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_63_buf (.a(edt_scan_in_buf_in[63]),
                                                                 .o(edt_scan_in[63]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_64_buf (.a(edt_scan_in_buf_in[64]),
                                                                 .o(edt_scan_in[64]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_65_buf (.a(edt_scan_in_buf_in[65]),
                                                                 .o(edt_scan_in[65]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_66_buf (.a(edt_scan_in_buf_in[66]),
                                                                 .o(edt_scan_in[66]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_67_buf (.a(edt_scan_in_buf_in[67]),
                                                                 .o(edt_scan_in[67]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_68_buf (.a(edt_scan_in_buf_in[68]),
                                                                 .o(edt_scan_in[68]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_69_buf (.a(edt_scan_in_buf_in[69]),
                                                                 .o(edt_scan_in[69]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_70_buf (.a(edt_scan_in_buf_in[70]),
                                                                 .o(edt_scan_in[70]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_71_buf (.a(edt_scan_in_buf_in[71]),
                                                                 .o(edt_scan_in[71]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_72_buf (.a(edt_scan_in_buf_in[72]),
                                                                 .o(edt_scan_in[72]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_73_buf (.a(edt_scan_in_buf_in[73]),
                                                                 .o(edt_scan_in[73]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_74_buf (.a(edt_scan_in_buf_in[74]),
                                                                 .o(edt_scan_in[74]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_75_buf (.a(edt_scan_in_buf_in[75]),
                                                                 .o(edt_scan_in[75]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_76_buf (.a(edt_scan_in_buf_in[76]),
                                                                 .o(edt_scan_in[76]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_77_buf (.a(edt_scan_in_buf_in[77]),
                                                                 .o(edt_scan_in[77]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_78_buf (.a(edt_scan_in_buf_in[78]),
                                                                 .o(edt_scan_in[78]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_79_buf (.a(edt_scan_in_buf_in[79]),
                                                                 .o(edt_scan_in[79]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_80_buf (.a(edt_scan_in_buf_in[80]),
                                                                 .o(edt_scan_in[80]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_81_buf (.a(edt_scan_in_buf_in[81]),
                                                                 .o(edt_scan_in[81]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_82_buf (.a(edt_scan_in_buf_in[82]),
                                                                 .o(edt_scan_in[82]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_83_buf (.a(edt_scan_in_buf_in[83]),
                                                                 .o(edt_scan_in[83]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_84_buf (.a(edt_scan_in_buf_in[84]),
                                                                 .o(edt_scan_in[84]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_85_buf (.a(edt_scan_in_buf_in[85]),
                                                                 .o(edt_scan_in[85]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_86_buf (.a(edt_scan_in_buf_in[86]),
                                                                 .o(edt_scan_in[86]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_87_buf (.a(edt_scan_in_buf_in[87]),
                                                                 .o(edt_scan_in[87]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_88_buf (.a(edt_scan_in_buf_in[88]),
                                                                 .o(edt_scan_in[88]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_89_buf (.a(edt_scan_in_buf_in[89]),
                                                                 .o(edt_scan_in[89]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_90_buf (.a(edt_scan_in_buf_in[90]),
                                                                 .o(edt_scan_in[90]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_91_buf (.a(edt_scan_in_buf_in[91]),
                                                                 .o(edt_scan_in[91]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_92_buf (.a(edt_scan_in_buf_in[92]),
                                                                 .o(edt_scan_in[92]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_93_buf (.a(edt_scan_in_buf_in[93]),
                                                                 .o(edt_scan_in[93]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_94_buf (.a(edt_scan_in_buf_in[94]),
                                                                 .o(edt_scan_in[94]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_95_buf (.a(edt_scan_in_buf_in[95]),
                                                                 .o(edt_scan_in[95]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_96_buf (.a(edt_scan_in_buf_in[96]),
                                                                 .o(edt_scan_in[96]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_97_buf (.a(edt_scan_in_buf_in[97]),
                                                                 .o(edt_scan_in[97]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_98_buf (.a(edt_scan_in_buf_in[98]),
                                                                 .o(edt_scan_in[98]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_99_buf (.a(edt_scan_in_buf_in[99]),
                                                                 .o(edt_scan_in[99]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_100_buf (.a(edt_scan_in_buf_in[100]),
                                                                  .o(edt_scan_in[100]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_101_buf (.a(edt_scan_in_buf_in[101]),
                                                                  .o(edt_scan_in[101]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_102_buf (.a(edt_scan_in_buf_in[102]),
                                                                  .o(edt_scan_in[102]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_103_buf (.a(edt_scan_in_buf_in[103]),
                                                                  .o(edt_scan_in[103]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_104_buf (.a(edt_scan_in_buf_in[104]),
                                                                  .o(edt_scan_in[104]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_105_buf (.a(edt_scan_in_buf_in[105]),
                                                                  .o(edt_scan_in[105]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_106_buf (.a(edt_scan_in_buf_in[106]),
                                                                  .o(edt_scan_in[106]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_107_buf (.a(edt_scan_in_buf_in[107]),
                                                                  .o(edt_scan_in[107]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_108_buf (.a(edt_scan_in_buf_in[108]),
                                                                  .o(edt_scan_in[108]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_109_buf (.a(edt_scan_in_buf_in[109]),
                                                                  .o(edt_scan_in[109]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_110_buf (.a(edt_scan_in_buf_in[110]),
                                                                  .o(edt_scan_in[110]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_111_buf (.a(edt_scan_in_buf_in[111]),
                                                                  .o(edt_scan_in[111]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_112_buf (.a(edt_scan_in_buf_in[112]),
                                                                  .o(edt_scan_in[112]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_113_buf (.a(edt_scan_in_buf_in[113]),
                                                                  .o(edt_scan_in[113]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_114_buf (.a(edt_scan_in_buf_in[114]),
                                                                  .o(edt_scan_in[114]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_115_buf (.a(edt_scan_in_buf_in[115]),
                                                                  .o(edt_scan_in[115]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_116_buf (.a(edt_scan_in_buf_in[116]),
                                                                  .o(edt_scan_in[116]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_117_buf (.a(edt_scan_in_buf_in[117]),
                                                                  .o(edt_scan_in[117]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_118_buf (.a(edt_scan_in_buf_in[118]),
                                                                  .o(edt_scan_in[118]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_119_buf (.a(edt_scan_in_buf_in[119]),
                                                                  .o(edt_scan_in[119]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_120_buf (.a(edt_scan_in_buf_in[120]),
                                                                  .o(edt_scan_in[120]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_121_buf (.a(edt_scan_in_buf_in[121]),
                                                                  .o(edt_scan_in[121]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_122_buf (.a(edt_scan_in_buf_in[122]),
                                                                  .o(edt_scan_in[122]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_123_buf (.a(edt_scan_in_buf_in[123]),
                                                                  .o(edt_scan_in[123]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_124_buf (.a(edt_scan_in_buf_in[124]),
                                                                  .o(edt_scan_in[124]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_125_buf (.a(edt_scan_in_buf_in[125]),
                                                                  .o(edt_scan_in[125]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_126_buf (.a(edt_scan_in_buf_in[126]),
                                                                  .o(edt_scan_in[126]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_127_buf (.a(edt_scan_in_buf_in[127]),
                                                                  .o(edt_scan_in[127]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_128_buf (.a(edt_scan_in_buf_in[128]),
                                                                  .o(edt_scan_in[128]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_129_buf (.a(edt_scan_in_buf_in[129]),
                                                                  .o(edt_scan_in[129]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_130_buf (.a(edt_scan_in_buf_in[130]),
                                                                  .o(edt_scan_in[130]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_131_buf (.a(edt_scan_in_buf_in[131]),
                                                                  .o(edt_scan_in[131]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_132_buf (.a(edt_scan_in_buf_in[132]),
                                                                  .o(edt_scan_in[132]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_133_buf (.a(edt_scan_in_buf_in[133]),
                                                                  .o(edt_scan_in[133]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_134_buf (.a(edt_scan_in_buf_in[134]),
                                                                  .o(edt_scan_in[134]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_135_buf (.a(edt_scan_in_buf_in[135]),
                                                                  .o(edt_scan_in[135]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_136_buf (.a(edt_scan_in_buf_in[136]),
                                                                  .o(edt_scan_in[136]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_137_buf (.a(edt_scan_in_buf_in[137]),
                                                                  .o(edt_scan_in[137]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_138_buf (.a(edt_scan_in_buf_in[138]),
                                                                  .o(edt_scan_in[138]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_139_buf (.a(edt_scan_in_buf_in[139]),
                                                                  .o(edt_scan_in[139]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_140_buf (.a(edt_scan_in_buf_in[140]),
                                                                  .o(edt_scan_in[140]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_141_buf (.a(edt_scan_in_buf_in[141]),
                                                                  .o(edt_scan_in[141]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_142_buf (.a(edt_scan_in_buf_in[142]),
                                                                  .o(edt_scan_in[142]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_143_buf (.a(edt_scan_in_buf_in[143]),
                                                                  .o(edt_scan_in[143]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_144_buf (.a(edt_scan_in_buf_in[144]),
                                                                  .o(edt_scan_in[144]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_145_buf (.a(edt_scan_in_buf_in[145]),
                                                                  .o(edt_scan_in[145]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_146_buf (.a(edt_scan_in_buf_in[146]),
                                                                  .o(edt_scan_in[146]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_147_buf (.a(edt_scan_in_buf_in[147]),
                                                                  .o(edt_scan_in[147]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_148_buf (.a(edt_scan_in_buf_in[148]),
                                                                  .o(edt_scan_in[148]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_149_buf (.a(edt_scan_in_buf_in[149]),
                                                                  .o(edt_scan_in[149]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_150_buf (.a(edt_scan_in_buf_in[150]),
                                                                  .o(edt_scan_in[150]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_151_buf (.a(edt_scan_in_buf_in[151]),
                                                                  .o(edt_scan_in[151]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_152_buf (.a(edt_scan_in_buf_in[152]),
                                                                  .o(edt_scan_in[152]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_153_buf (.a(edt_scan_in_buf_in[153]),
                                                                  .o(edt_scan_in[153]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_154_buf (.a(edt_scan_in_buf_in[154]),
                                                                  .o(edt_scan_in[154]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_155_buf (.a(edt_scan_in_buf_in[155]),
                                                                  .o(edt_scan_in[155]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_156_buf (.a(edt_scan_in_buf_in[156]),
                                                                  .o(edt_scan_in[156]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_157_buf (.a(edt_scan_in_buf_in[157]),
                                                                  .o(edt_scan_in[157]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_158_buf (.a(edt_scan_in_buf_in[158]),
                                                                  .o(edt_scan_in[158]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_159_buf (.a(edt_scan_in_buf_in[159]),
                                                                  .o(edt_scan_in[159]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_160_buf (.a(edt_scan_in_buf_in[160]),
                                                                  .o(edt_scan_in[160]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_161_buf (.a(edt_scan_in_buf_in[161]),
                                                                  .o(edt_scan_in[161]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_162_buf (.a(edt_scan_in_buf_in[162]),
                                                                  .o(edt_scan_in[162]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_163_buf (.a(edt_scan_in_buf_in[163]),
                                                                  .o(edt_scan_in[163]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_164_buf (.a(edt_scan_in_buf_in[164]),
                                                                  .o(edt_scan_in[164]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_165_buf (.a(edt_scan_in_buf_in[165]),
                                                                  .o(edt_scan_in[165]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_166_buf (.a(edt_scan_in_buf_in[166]),
                                                                  .o(edt_scan_in[166]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_167_buf (.a(edt_scan_in_buf_in[167]),
                                                                  .o(edt_scan_in[167]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_168_buf (.a(edt_scan_in_buf_in[168]),
                                                                  .o(edt_scan_in[168]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_169_buf (.a(edt_scan_in_buf_in[169]),
                                                                  .o(edt_scan_in[169]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_170_buf (.a(edt_scan_in_buf_in[170]),
                                                                  .o(edt_scan_in[170]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_171_buf (.a(edt_scan_in_buf_in[171]),
                                                                  .o(edt_scan_in[171]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_172_buf (.a(edt_scan_in_buf_in[172]),
                                                                  .o(edt_scan_in[172]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_173_buf (.a(edt_scan_in_buf_in[173]),
                                                                  .o(edt_scan_in[173]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_174_buf (.a(edt_scan_in_buf_in[174]),
                                                                  .o(edt_scan_in[174]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_175_buf (.a(edt_scan_in_buf_in[175]),
                                                                  .o(edt_scan_in[175]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_176_buf (.a(edt_scan_in_buf_in[176]),
                                                                  .o(edt_scan_in[176]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_177_buf (.a(edt_scan_in_buf_in[177]),
                                                                  .o(edt_scan_in[177]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_178_buf (.a(edt_scan_in_buf_in[178]),
                                                                  .o(edt_scan_in[178]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_179_buf (.a(edt_scan_in_buf_in[179]),
                                                                  .o(edt_scan_in[179]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_180_buf (.a(edt_scan_in_buf_in[180]),
                                                                  .o(edt_scan_in[180]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_181_buf (.a(edt_scan_in_buf_in[181]),
                                                                  .o(edt_scan_in[181]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_182_buf (.a(edt_scan_in_buf_in[182]),
                                                                  .o(edt_scan_in[182]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_183_buf (.a(edt_scan_in_buf_in[183]),
                                                                  .o(edt_scan_in[183]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_184_buf (.a(edt_scan_in_buf_in[184]),
                                                                  .o(edt_scan_in[184]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_185_buf (.a(edt_scan_in_buf_in[185]),
                                                                  .o(edt_scan_in[185]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_186_buf (.a(edt_scan_in_buf_in[186]),
                                                                  .o(edt_scan_in[186]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_187_buf (.a(edt_scan_in_buf_in[187]),
                                                                  .o(edt_scan_in[187]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_188_buf (.a(edt_scan_in_buf_in[188]),
                                                                  .o(edt_scan_in[188]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_189_buf (.a(edt_scan_in_buf_in[189]),
                                                                  .o(edt_scan_in[189]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_190_buf (.a(edt_scan_in_buf_in[190]),
                                                                  .o(edt_scan_in[190]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_191_buf (.a(edt_scan_in_buf_in[191]),
                                                                  .o(edt_scan_in[191]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_192_buf (.a(edt_scan_in_buf_in[192]),
                                                                  .o(edt_scan_in[192]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_193_buf (.a(edt_scan_in_buf_in[193]),
                                                                  .o(edt_scan_in[193]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_194_buf (.a(edt_scan_in_buf_in[194]),
                                                                  .o(edt_scan_in[194]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_195_buf (.a(edt_scan_in_buf_in[195]),
                                                                  .o(edt_scan_in[195]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_196_buf (.a(edt_scan_in_buf_in[196]),
                                                                  .o(edt_scan_in[196]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_197_buf (.a(edt_scan_in_buf_in[197]),
                                                                  .o(edt_scan_in[197]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_198_buf (.a(edt_scan_in_buf_in[198]),
                                                                  .o(edt_scan_in[198]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_199_buf (.a(edt_scan_in_buf_in[199]),
                                                                  .o(edt_scan_in[199]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_200_buf (.a(edt_scan_in_buf_in[200]),
                                                                  .o(edt_scan_in[200]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_201_buf (.a(edt_scan_in_buf_in[201]),
                                                                  .o(edt_scan_in[201]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_202_buf (.a(edt_scan_in_buf_in[202]),
                                                                  .o(edt_scan_in[202]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_203_buf (.a(edt_scan_in_buf_in[203]),
                                                                  .o(edt_scan_in[203]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_204_buf (.a(edt_scan_in_buf_in[204]),
                                                                  .o(edt_scan_in[204]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_205_buf (.a(edt_scan_in_buf_in[205]),
                                                                  .o(edt_scan_in[205]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_206_buf (.a(edt_scan_in_buf_in[206]),
                                                                  .o(edt_scan_in[206]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_207_buf (.a(edt_scan_in_buf_in[207]),
                                                                  .o(edt_scan_in[207]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_208_buf (.a(edt_scan_in_buf_in[208]),
                                                                  .o(edt_scan_in[208]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_209_buf (.a(edt_scan_in_buf_in[209]),
                                                                  .o(edt_scan_in[209]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_210_buf (.a(edt_scan_in_buf_in[210]),
                                                                  .o(edt_scan_in[210]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_211_buf (.a(edt_scan_in_buf_in[211]),
                                                                  .o(edt_scan_in[211]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_212_buf (.a(edt_scan_in_buf_in[212]),
                                                                  .o(edt_scan_in[212]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_213_buf (.a(edt_scan_in_buf_in[213]),
                                                                  .o(edt_scan_in[213]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_214_buf (.a(edt_scan_in_buf_in[214]),
                                                                  .o(edt_scan_in[214]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_215_buf (.a(edt_scan_in_buf_in[215]),
                                                                  .o(edt_scan_in[215]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_216_buf (.a(edt_scan_in_buf_in[216]),
                                                                  .o(edt_scan_in[216]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_217_buf (.a(edt_scan_in_buf_in[217]),
                                                                  .o(edt_scan_in[217]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_218_buf (.a(edt_scan_in_buf_in[218]),
                                                                  .o(edt_scan_in[218]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_219_buf (.a(edt_scan_in_buf_in[219]),
                                                                  .o(edt_scan_in[219]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_220_buf (.a(edt_scan_in_buf_in[220]),
                                                                  .o(edt_scan_in[220]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_221_buf (.a(edt_scan_in_buf_in[221]),
                                                                  .o(edt_scan_in[221]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_222_buf (.a(edt_scan_in_buf_in[222]),
                                                                  .o(edt_scan_in[222]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_223_buf (.a(edt_scan_in_buf_in[223]),
                                                                  .o(edt_scan_in[223]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_224_buf (.a(edt_scan_in_buf_in[224]),
                                                                  .o(edt_scan_in[224]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_225_buf (.a(edt_scan_in_buf_in[225]),
                                                                  .o(edt_scan_in[225]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_226_buf (.a(edt_scan_in_buf_in[226]),
                                                                  .o(edt_scan_in[226]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_227_buf (.a(edt_scan_in_buf_in[227]),
                                                                  .o(edt_scan_in[227]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_228_buf (.a(edt_scan_in_buf_in[228]),
                                                                  .o(edt_scan_in[228]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_229_buf (.a(edt_scan_in_buf_in[229]),
                                                                  .o(edt_scan_in[229]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_230_buf (.a(edt_scan_in_buf_in[230]),
                                                                  .o(edt_scan_in[230]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_231_buf (.a(edt_scan_in_buf_in[231]),
                                                                  .o(edt_scan_in[231]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_232_buf (.a(edt_scan_in_buf_in[232]),
                                                                  .o(edt_scan_in[232]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_233_buf (.a(edt_scan_in_buf_in[233]),
                                                                  .o(edt_scan_in[233]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_234_buf (.a(edt_scan_in_buf_in[234]),
                                                                  .o(edt_scan_in[234]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_235_buf (.a(edt_scan_in_buf_in[235]),
                                                                  .o(edt_scan_in[235]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_236_buf (.a(edt_scan_in_buf_in[236]),
                                                                  .o(edt_scan_in[236]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_237_buf (.a(edt_scan_in_buf_in[237]),
                                                                  .o(edt_scan_in[237]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_238_buf (.a(edt_scan_in_buf_in[238]),
                                                                  .o(edt_scan_in[238]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_239_buf (.a(edt_scan_in_buf_in[239]),
                                                                  .o(edt_scan_in[239]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_240_buf (.a(edt_scan_in_buf_in[240]),
                                                                  .o(edt_scan_in[240]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_241_buf (.a(edt_scan_in_buf_in[241]),
                                                                  .o(edt_scan_in[241]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_242_buf (.a(edt_scan_in_buf_in[242]),
                                                                  .o(edt_scan_in[242]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_243_buf (.a(edt_scan_in_buf_in[243]),
                                                                  .o(edt_scan_in[243]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_244_buf (.a(edt_scan_in_buf_in[244]),
                                                                  .o(edt_scan_in[244]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_245_buf (.a(edt_scan_in_buf_in[245]),
                                                                  .o(edt_scan_in[245]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_246_buf (.a(edt_scan_in_buf_in[246]),
                                                                  .o(edt_scan_in[246]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_247_buf (.a(edt_scan_in_buf_in[247]),
                                                                  .o(edt_scan_in[247]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_248_buf (.a(edt_scan_in_buf_in[248]),
                                                                  .o(edt_scan_in[248]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_249_buf (.a(edt_scan_in_buf_in[249]),
                                                                  .o(edt_scan_in[249]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_250_buf (.a(edt_scan_in_buf_in[250]),
                                                                  .o(edt_scan_in[250]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_251_buf (.a(edt_scan_in_buf_in[251]),
                                                                  .o(edt_scan_in[251]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_252_buf (.a(edt_scan_in_buf_in[252]),
                                                                  .o(edt_scan_in[252]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_253_buf (.a(edt_scan_in_buf_in[253]),
                                                                  .o(edt_scan_in[253]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_254_buf (.a(edt_scan_in_buf_in[254]),
                                                                  .o(edt_scan_in[254]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_255_buf (.a(edt_scan_in_buf_in[255]),
                                                                  .o(edt_scan_in[255]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_256_buf (.a(edt_scan_in_buf_in[256]),
                                                                  .o(edt_scan_in[256]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_257_buf (.a(edt_scan_in_buf_in[257]),
                                                                  .o(edt_scan_in[257]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_258_buf (.a(edt_scan_in_buf_in[258]),
                                                                  .o(edt_scan_in[258]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_259_buf (.a(edt_scan_in_buf_in[259]),
                                                                  .o(edt_scan_in[259]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_260_buf (.a(edt_scan_in_buf_in[260]),
                                                                  .o(edt_scan_in[260]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_261_buf (.a(edt_scan_in_buf_in[261]),
                                                                  .o(edt_scan_in[261]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_262_buf (.a(edt_scan_in_buf_in[262]),
                                                                  .o(edt_scan_in[262]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_263_buf (.a(edt_scan_in_buf_in[263]),
                                                                  .o(edt_scan_in[263]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_264_buf (.a(edt_scan_in_buf_in[264]),
                                                                  .o(edt_scan_in[264]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_265_buf (.a(edt_scan_in_buf_in[265]),
                                                                  .o(edt_scan_in[265]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_266_buf (.a(edt_scan_in_buf_in[266]),
                                                                  .o(edt_scan_in[266]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_267_buf (.a(edt_scan_in_buf_in[267]),
                                                                  .o(edt_scan_in[267]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_268_buf (.a(edt_scan_in_buf_in[268]),
                                                                  .o(edt_scan_in[268]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_269_buf (.a(edt_scan_in_buf_in[269]),
                                                                  .o(edt_scan_in[269]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_270_buf (.a(edt_scan_in_buf_in[270]),
                                                                  .o(edt_scan_in[270]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_271_buf (.a(edt_scan_in_buf_in[271]),
                                                                  .o(edt_scan_in[271]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_272_buf (.a(edt_scan_in_buf_in[272]),
                                                                  .o(edt_scan_in[272]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_273_buf (.a(edt_scan_in_buf_in[273]),
                                                                  .o(edt_scan_in[273]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_274_buf (.a(edt_scan_in_buf_in[274]),
                                                                  .o(edt_scan_in[274]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_275_buf (.a(edt_scan_in_buf_in[275]),
                                                                  .o(edt_scan_in[275]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_276_buf (.a(edt_scan_in_buf_in[276]),
                                                                  .o(edt_scan_in[276]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_277_buf (.a(edt_scan_in_buf_in[277]),
                                                                  .o(edt_scan_in[277]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_278_buf (.a(edt_scan_in_buf_in[278]),
                                                                  .o(edt_scan_in[278]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_279_buf (.a(edt_scan_in_buf_in[279]),
                                                                  .o(edt_scan_in[279]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_280_buf (.a(edt_scan_in_buf_in[280]),
                                                                  .o(edt_scan_in[280]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_281_buf (.a(edt_scan_in_buf_in[281]),
                                                                  .o(edt_scan_in[281]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_282_buf (.a(edt_scan_in_buf_in[282]),
                                                                  .o(edt_scan_in[282]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_283_buf (.a(edt_scan_in_buf_in[283]),
                                                                  .o(edt_scan_in[283]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_284_buf (.a(edt_scan_in_buf_in[284]),
                                                                  .o(edt_scan_in[284]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_285_buf (.a(edt_scan_in_buf_in[285]),
                                                                  .o(edt_scan_in[285]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_286_buf (.a(edt_scan_in_buf_in[286]),
                                                                  .o(edt_scan_in[286]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_287_buf (.a(edt_scan_in_buf_in[287]),
                                                                  .o(edt_scan_in[287]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_288_buf (.a(edt_scan_in_buf_in[288]),
                                                                  .o(edt_scan_in[288]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_289_buf (.a(edt_scan_in_buf_in[289]),
                                                                  .o(edt_scan_in[289]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_290_buf (.a(edt_scan_in_buf_in[290]),
                                                                  .o(edt_scan_in[290]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_291_buf (.a(edt_scan_in_buf_in[291]),
                                                                  .o(edt_scan_in[291]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_292_buf (.a(edt_scan_in_buf_in[292]),
                                                                  .o(edt_scan_in[292]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_293_buf (.a(edt_scan_in_buf_in[293]),
                                                                  .o(edt_scan_in[293]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_294_buf (.a(edt_scan_in_buf_in[294]),
                                                                  .o(edt_scan_in[294]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_295_buf (.a(edt_scan_in_buf_in[295]),
                                                                  .o(edt_scan_in[295]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_296_buf (.a(edt_scan_in_buf_in[296]),
                                                                  .o(edt_scan_in[296]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_297_buf (.a(edt_scan_in_buf_in[297]),
                                                                  .o(edt_scan_in[297]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_298_buf (.a(edt_scan_in_buf_in[298]),
                                                                  .o(edt_scan_in[298]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_299_buf (.a(edt_scan_in_buf_in[299]),
                                                                  .o(edt_scan_in[299]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_300_buf (.a(edt_scan_in_buf_in[300]),
                                                                  .o(edt_scan_in[300]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_301_buf (.a(edt_scan_in_buf_in[301]),
                                                                  .o(edt_scan_in[301]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_302_buf (.a(edt_scan_in_buf_in[302]),
                                                                  .o(edt_scan_in[302]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_303_buf (.a(edt_scan_in_buf_in[303]),
                                                                  .o(edt_scan_in[303]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_304_buf (.a(edt_scan_in_buf_in[304]),
                                                                  .o(edt_scan_in[304]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_305_buf (.a(edt_scan_in_buf_in[305]),
                                                                  .o(edt_scan_in[305]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_306_buf (.a(edt_scan_in_buf_in[306]),
                                                                  .o(edt_scan_in[306]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_307_buf (.a(edt_scan_in_buf_in[307]),
                                                                  .o(edt_scan_in[307]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_308_buf (.a(edt_scan_in_buf_in[308]),
                                                                  .o(edt_scan_in[308]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_309_buf (.a(edt_scan_in_buf_in[309]),
                                                                  .o(edt_scan_in[309]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_310_buf (.a(edt_scan_in_buf_in[310]),
                                                                  .o(edt_scan_in[310]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_311_buf (.a(edt_scan_in_buf_in[311]),
                                                                  .o(edt_scan_in[311]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_312_buf (.a(edt_scan_in_buf_in[312]),
                                                                  .o(edt_scan_in[312]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_313_buf (.a(edt_scan_in_buf_in[313]),
                                                                  .o(edt_scan_in[313]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_314_buf (.a(edt_scan_in_buf_in[314]),
                                                                  .o(edt_scan_in[314]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_315_buf (.a(edt_scan_in_buf_in[315]),
                                                                  .o(edt_scan_in[315]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_316_buf (.a(edt_scan_in_buf_in[316]),
                                                                  .o(edt_scan_in[316]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_317_buf (.a(edt_scan_in_buf_in[317]),
                                                                  .o(edt_scan_in[317]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_318_buf (.a(edt_scan_in_buf_in[318]),
                                                                  .o(edt_scan_in[318]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_319_buf (.a(edt_scan_in_buf_in[319]),
                                                                  .o(edt_scan_in[319]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_320_buf (.a(edt_scan_in_buf_in[320]),
                                                                  .o(edt_scan_in[320]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_321_buf (.a(edt_scan_in_buf_in[321]),
                                                                  .o(edt_scan_in[321]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_322_buf (.a(edt_scan_in_buf_in[322]),
                                                                  .o(edt_scan_in[322]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_323_buf (.a(edt_scan_in_buf_in[323]),
                                                                  .o(edt_scan_in[323]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_324_buf (.a(edt_scan_in_buf_in[324]),
                                                                  .o(edt_scan_in[324]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_325_buf (.a(edt_scan_in_buf_in[325]),
                                                                  .o(edt_scan_in[325]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_326_buf (.a(edt_scan_in_buf_in[326]),
                                                                  .o(edt_scan_in[326]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_327_buf (.a(edt_scan_in_buf_in[327]),
                                                                  .o(edt_scan_in[327]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_328_buf (.a(edt_scan_in_buf_in[328]),
                                                                  .o(edt_scan_in[328]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_329_buf (.a(edt_scan_in_buf_in[329]),
                                                                  .o(edt_scan_in[329]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_330_buf (.a(edt_scan_in_buf_in[330]),
                                                                  .o(edt_scan_in[330]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_331_buf (.a(edt_scan_in_buf_in[331]),
                                                                  .o(edt_scan_in[331]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_332_buf (.a(edt_scan_in_buf_in[332]),
                                                                  .o(edt_scan_in[332]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_333_buf (.a(edt_scan_in_buf_in[333]),
                                                                  .o(edt_scan_in[333]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_334_buf (.a(edt_scan_in_buf_in[334]),
                                                                  .o(edt_scan_in[334]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_335_buf (.a(edt_scan_in_buf_in[335]),
                                                                  .o(edt_scan_in[335]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_336_buf (.a(edt_scan_in_buf_in[336]),
                                                                  .o(edt_scan_in[336]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_337_buf (.a(edt_scan_in_buf_in[337]),
                                                                  .o(edt_scan_in[337]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_338_buf (.a(edt_scan_in_buf_in[338]),
                                                                  .o(edt_scan_in[338]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_339_buf (.a(edt_scan_in_buf_in[339]),
                                                                  .o(edt_scan_in[339]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_340_buf (.a(edt_scan_in_buf_in[340]),
                                                                  .o(edt_scan_in[340]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_341_buf (.a(edt_scan_in_buf_in[341]),
                                                                  .o(edt_scan_in[341]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_342_buf (.a(edt_scan_in_buf_in[342]),
                                                                  .o(edt_scan_in[342]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_343_buf (.a(edt_scan_in_buf_in[343]),
                                                                  .o(edt_scan_in[343]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_344_buf (.a(edt_scan_in_buf_in[344]),
                                                                  .o(edt_scan_in[344]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_345_buf (.a(edt_scan_in_buf_in[345]),
                                                                  .o(edt_scan_in[345]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_346_buf (.a(edt_scan_in_buf_in[346]),
                                                                  .o(edt_scan_in[346]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_347_buf (.a(edt_scan_in_buf_in[347]),
                                                                  .o(edt_scan_in[347]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_348_buf (.a(edt_scan_in_buf_in[348]),
                                                                  .o(edt_scan_in[348]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_349_buf (.a(edt_scan_in_buf_in[349]),
                                                                  .o(edt_scan_in[349]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_350_buf (.a(edt_scan_in_buf_in[350]),
                                                                  .o(edt_scan_in[350]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_351_buf (.a(edt_scan_in_buf_in[351]),
                                                                  .o(edt_scan_in[351]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_352_buf (.a(edt_scan_in_buf_in[352]),
                                                                  .o(edt_scan_in[352]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_353_buf (.a(edt_scan_in_buf_in[353]),
                                                                  .o(edt_scan_in[353]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_354_buf (.a(edt_scan_in_buf_in[354]),
                                                                  .o(edt_scan_in[354]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_355_buf (.a(edt_scan_in_buf_in[355]),
                                                                  .o(edt_scan_in[355]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_356_buf (.a(edt_scan_in_buf_in[356]),
                                                                  .o(edt_scan_in[356]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_357_buf (.a(edt_scan_in_buf_in[357]),
                                                                  .o(edt_scan_in[357]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_358_buf (.a(edt_scan_in_buf_in[358]),
                                                                  .o(edt_scan_in[358]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_359_buf (.a(edt_scan_in_buf_in[359]),
                                                                  .o(edt_scan_in[359]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_360_buf (.a(edt_scan_in_buf_in[360]),
                                                                  .o(edt_scan_in[360]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_361_buf (.a(edt_scan_in_buf_in[361]),
                                                                  .o(edt_scan_in[361]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_362_buf (.a(edt_scan_in_buf_in[362]),
                                                                  .o(edt_scan_in[362]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_363_buf (.a(edt_scan_in_buf_in[363]),
                                                                  .o(edt_scan_in[363]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_364_buf (.a(edt_scan_in_buf_in[364]),
                                                                  .o(edt_scan_in[364]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_365_buf (.a(edt_scan_in_buf_in[365]),
                                                                  .o(edt_scan_in[365]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_366_buf (.a(edt_scan_in_buf_in[366]),
                                                                  .o(edt_scan_in[366]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_367_buf (.a(edt_scan_in_buf_in[367]),
                                                                  .o(edt_scan_in[367]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_368_buf (.a(edt_scan_in_buf_in[368]),
                                                                  .o(edt_scan_in[368]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_369_buf (.a(edt_scan_in_buf_in[369]),
                                                                  .o(edt_scan_in[369]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_in_370_buf (.a(edt_scan_in_buf_in[370]),
                                                                  .o(edt_scan_in[370]));

   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_0_buf (.a(edt_scan_out[0]),
                                                                 .o(edt_scan_out_buf_out[0]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_1_buf (.a(edt_scan_out[1]),
                                                                 .o(edt_scan_out_buf_out[1]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_2_buf (.a(edt_scan_out[2]),
                                                                 .o(edt_scan_out_buf_out[2]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_3_buf (.a(edt_scan_out[3]),
                                                                 .o(edt_scan_out_buf_out[3]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_4_buf (.a(edt_scan_out[4]),
                                                                 .o(edt_scan_out_buf_out[4]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_5_buf (.a(edt_scan_out[5]),
                                                                 .o(edt_scan_out_buf_out[5]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_6_buf (.a(edt_scan_out[6]),
                                                                 .o(edt_scan_out_buf_out[6]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_7_buf (.a(edt_scan_out[7]),
                                                                 .o(edt_scan_out_buf_out[7]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_8_buf (.a(edt_scan_out[8]),
                                                                 .o(edt_scan_out_buf_out[8]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_9_buf (.a(edt_scan_out[9]),
                                                                 .o(edt_scan_out_buf_out[9]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_10_buf (.a(edt_scan_out[10]),
                                                                  .o(edt_scan_out_buf_out[10]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_11_buf (.a(edt_scan_out[11]),
                                                                  .o(edt_scan_out_buf_out[11]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_12_buf (.a(edt_scan_out[12]),
                                                                  .o(edt_scan_out_buf_out[12]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_13_buf (.a(edt_scan_out[13]),
                                                                  .o(edt_scan_out_buf_out[13]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_14_buf (.a(edt_scan_out[14]),
                                                                  .o(edt_scan_out_buf_out[14]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_15_buf (.a(edt_scan_out[15]),
                                                                  .o(edt_scan_out_buf_out[15]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_16_buf (.a(edt_scan_out[16]),
                                                                  .o(edt_scan_out_buf_out[16]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_17_buf (.a(edt_scan_out[17]),
                                                                  .o(edt_scan_out_buf_out[17]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_18_buf (.a(edt_scan_out[18]),
                                                                  .o(edt_scan_out_buf_out[18]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_19_buf (.a(edt_scan_out[19]),
                                                                  .o(edt_scan_out_buf_out[19]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_20_buf (.a(edt_scan_out[20]),
                                                                  .o(edt_scan_out_buf_out[20]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_21_buf (.a(edt_scan_out[21]),
                                                                  .o(edt_scan_out_buf_out[21]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_22_buf (.a(edt_scan_out[22]),
                                                                  .o(edt_scan_out_buf_out[22]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_23_buf (.a(edt_scan_out[23]),
                                                                  .o(edt_scan_out_buf_out[23]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_24_buf (.a(edt_scan_out[24]),
                                                                  .o(edt_scan_out_buf_out[24]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_25_buf (.a(edt_scan_out[25]),
                                                                  .o(edt_scan_out_buf_out[25]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_26_buf (.a(edt_scan_out[26]),
                                                                  .o(edt_scan_out_buf_out[26]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_27_buf (.a(edt_scan_out[27]),
                                                                  .o(edt_scan_out_buf_out[27]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_28_buf (.a(edt_scan_out[28]),
                                                                  .o(edt_scan_out_buf_out[28]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_29_buf (.a(edt_scan_out[29]),
                                                                  .o(edt_scan_out_buf_out[29]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_30_buf (.a(edt_scan_out[30]),
                                                                  .o(edt_scan_out_buf_out[30]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_31_buf (.a(edt_scan_out[31]),
                                                                  .o(edt_scan_out_buf_out[31]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_32_buf (.a(edt_scan_out[32]),
                                                                  .o(edt_scan_out_buf_out[32]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_33_buf (.a(edt_scan_out[33]),
                                                                  .o(edt_scan_out_buf_out[33]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_34_buf (.a(edt_scan_out[34]),
                                                                  .o(edt_scan_out_buf_out[34]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_35_buf (.a(edt_scan_out[35]),
                                                                  .o(edt_scan_out_buf_out[35]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_36_buf (.a(edt_scan_out[36]),
                                                                  .o(edt_scan_out_buf_out[36]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_37_buf (.a(edt_scan_out[37]),
                                                                  .o(edt_scan_out_buf_out[37]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_38_buf (.a(edt_scan_out[38]),
                                                                  .o(edt_scan_out_buf_out[38]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_39_buf (.a(edt_scan_out[39]),
                                                                  .o(edt_scan_out_buf_out[39]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_40_buf (.a(edt_scan_out[40]),
                                                                  .o(edt_scan_out_buf_out[40]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_41_buf (.a(edt_scan_out[41]),
                                                                  .o(edt_scan_out_buf_out[41]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_42_buf (.a(edt_scan_out[42]),
                                                                  .o(edt_scan_out_buf_out[42]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_43_buf (.a(edt_scan_out[43]),
                                                                  .o(edt_scan_out_buf_out[43]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_44_buf (.a(edt_scan_out[44]),
                                                                  .o(edt_scan_out_buf_out[44]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_45_buf (.a(edt_scan_out[45]),
                                                                  .o(edt_scan_out_buf_out[45]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_46_buf (.a(edt_scan_out[46]),
                                                                  .o(edt_scan_out_buf_out[46]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_47_buf (.a(edt_scan_out[47]),
                                                                  .o(edt_scan_out_buf_out[47]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_48_buf (.a(edt_scan_out[48]),
                                                                  .o(edt_scan_out_buf_out[48]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_49_buf (.a(edt_scan_out[49]),
                                                                  .o(edt_scan_out_buf_out[49]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_50_buf (.a(edt_scan_out[50]),
                                                                  .o(edt_scan_out_buf_out[50]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_51_buf (.a(edt_scan_out[51]),
                                                                  .o(edt_scan_out_buf_out[51]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_52_buf (.a(edt_scan_out[52]),
                                                                  .o(edt_scan_out_buf_out[52]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_53_buf (.a(edt_scan_out[53]),
                                                                  .o(edt_scan_out_buf_out[53]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_54_buf (.a(edt_scan_out[54]),
                                                                  .o(edt_scan_out_buf_out[54]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_55_buf (.a(edt_scan_out[55]),
                                                                  .o(edt_scan_out_buf_out[55]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_56_buf (.a(edt_scan_out[56]),
                                                                  .o(edt_scan_out_buf_out[56]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_57_buf (.a(edt_scan_out[57]),
                                                                  .o(edt_scan_out_buf_out[57]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_58_buf (.a(edt_scan_out[58]),
                                                                  .o(edt_scan_out_buf_out[58]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_59_buf (.a(edt_scan_out[59]),
                                                                  .o(edt_scan_out_buf_out[59]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_60_buf (.a(edt_scan_out[60]),
                                                                  .o(edt_scan_out_buf_out[60]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_61_buf (.a(edt_scan_out[61]),
                                                                  .o(edt_scan_out_buf_out[61]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_62_buf (.a(edt_scan_out[62]),
                                                                  .o(edt_scan_out_buf_out[62]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_63_buf (.a(edt_scan_out[63]),
                                                                  .o(edt_scan_out_buf_out[63]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_64_buf (.a(edt_scan_out[64]),
                                                                  .o(edt_scan_out_buf_out[64]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_65_buf (.a(edt_scan_out[65]),
                                                                  .o(edt_scan_out_buf_out[65]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_66_buf (.a(edt_scan_out[66]),
                                                                  .o(edt_scan_out_buf_out[66]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_67_buf (.a(edt_scan_out[67]),
                                                                  .o(edt_scan_out_buf_out[67]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_68_buf (.a(edt_scan_out[68]),
                                                                  .o(edt_scan_out_buf_out[68]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_69_buf (.a(edt_scan_out[69]),
                                                                  .o(edt_scan_out_buf_out[69]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_70_buf (.a(edt_scan_out[70]),
                                                                  .o(edt_scan_out_buf_out[70]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_71_buf (.a(edt_scan_out[71]),
                                                                  .o(edt_scan_out_buf_out[71]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_72_buf (.a(edt_scan_out[72]),
                                                                  .o(edt_scan_out_buf_out[72]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_73_buf (.a(edt_scan_out[73]),
                                                                  .o(edt_scan_out_buf_out[73]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_74_buf (.a(edt_scan_out[74]),
                                                                  .o(edt_scan_out_buf_out[74]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_75_buf (.a(edt_scan_out[75]),
                                                                  .o(edt_scan_out_buf_out[75]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_76_buf (.a(edt_scan_out[76]),
                                                                  .o(edt_scan_out_buf_out[76]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_77_buf (.a(edt_scan_out[77]),
                                                                  .o(edt_scan_out_buf_out[77]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_78_buf (.a(edt_scan_out[78]),
                                                                  .o(edt_scan_out_buf_out[78]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_79_buf (.a(edt_scan_out[79]),
                                                                  .o(edt_scan_out_buf_out[79]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_80_buf (.a(edt_scan_out[80]),
                                                                  .o(edt_scan_out_buf_out[80]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_81_buf (.a(edt_scan_out[81]),
                                                                  .o(edt_scan_out_buf_out[81]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_82_buf (.a(edt_scan_out[82]),
                                                                  .o(edt_scan_out_buf_out[82]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_83_buf (.a(edt_scan_out[83]),
                                                                  .o(edt_scan_out_buf_out[83]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_84_buf (.a(edt_scan_out[84]),
                                                                  .o(edt_scan_out_buf_out[84]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_85_buf (.a(edt_scan_out[85]),
                                                                  .o(edt_scan_out_buf_out[85]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_86_buf (.a(edt_scan_out[86]),
                                                                  .o(edt_scan_out_buf_out[86]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_87_buf (.a(edt_scan_out[87]),
                                                                  .o(edt_scan_out_buf_out[87]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_88_buf (.a(edt_scan_out[88]),
                                                                  .o(edt_scan_out_buf_out[88]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_89_buf (.a(edt_scan_out[89]),
                                                                  .o(edt_scan_out_buf_out[89]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_90_buf (.a(edt_scan_out[90]),
                                                                  .o(edt_scan_out_buf_out[90]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_91_buf (.a(edt_scan_out[91]),
                                                                  .o(edt_scan_out_buf_out[91]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_92_buf (.a(edt_scan_out[92]),
                                                                  .o(edt_scan_out_buf_out[92]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_93_buf (.a(edt_scan_out[93]),
                                                                  .o(edt_scan_out_buf_out[93]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_94_buf (.a(edt_scan_out[94]),
                                                                  .o(edt_scan_out_buf_out[94]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_95_buf (.a(edt_scan_out[95]),
                                                                  .o(edt_scan_out_buf_out[95]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_96_buf (.a(edt_scan_out[96]),
                                                                  .o(edt_scan_out_buf_out[96]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_97_buf (.a(edt_scan_out[97]),
                                                                  .o(edt_scan_out_buf_out[97]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_98_buf (.a(edt_scan_out[98]),
                                                                  .o(edt_scan_out_buf_out[98]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_99_buf (.a(edt_scan_out[99]),
                                                                  .o(edt_scan_out_buf_out[99]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_100_buf (.a(edt_scan_out[100]),
                                                                   .o(edt_scan_out_buf_out[100]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_101_buf (.a(edt_scan_out[101]),
                                                                   .o(edt_scan_out_buf_out[101]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_102_buf (.a(edt_scan_out[102]),
                                                                   .o(edt_scan_out_buf_out[102]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_103_buf (.a(edt_scan_out[103]),
                                                                   .o(edt_scan_out_buf_out[103]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_104_buf (.a(edt_scan_out[104]),
                                                                   .o(edt_scan_out_buf_out[104]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_105_buf (.a(edt_scan_out[105]),
                                                                   .o(edt_scan_out_buf_out[105]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_106_buf (.a(edt_scan_out[106]),
                                                                   .o(edt_scan_out_buf_out[106]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_107_buf (.a(edt_scan_out[107]),
                                                                   .o(edt_scan_out_buf_out[107]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_108_buf (.a(edt_scan_out[108]),
                                                                   .o(edt_scan_out_buf_out[108]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_109_buf (.a(edt_scan_out[109]),
                                                                   .o(edt_scan_out_buf_out[109]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_110_buf (.a(edt_scan_out[110]),
                                                                   .o(edt_scan_out_buf_out[110]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_111_buf (.a(edt_scan_out[111]),
                                                                   .o(edt_scan_out_buf_out[111]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_112_buf (.a(edt_scan_out[112]),
                                                                   .o(edt_scan_out_buf_out[112]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_113_buf (.a(edt_scan_out[113]),
                                                                   .o(edt_scan_out_buf_out[113]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_114_buf (.a(edt_scan_out[114]),
                                                                   .o(edt_scan_out_buf_out[114]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_115_buf (.a(edt_scan_out[115]),
                                                                   .o(edt_scan_out_buf_out[115]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_116_buf (.a(edt_scan_out[116]),
                                                                   .o(edt_scan_out_buf_out[116]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_117_buf (.a(edt_scan_out[117]),
                                                                   .o(edt_scan_out_buf_out[117]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_118_buf (.a(edt_scan_out[118]),
                                                                   .o(edt_scan_out_buf_out[118]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_119_buf (.a(edt_scan_out[119]),
                                                                   .o(edt_scan_out_buf_out[119]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_120_buf (.a(edt_scan_out[120]),
                                                                   .o(edt_scan_out_buf_out[120]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_121_buf (.a(edt_scan_out[121]),
                                                                   .o(edt_scan_out_buf_out[121]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_122_buf (.a(edt_scan_out[122]),
                                                                   .o(edt_scan_out_buf_out[122]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_123_buf (.a(edt_scan_out[123]),
                                                                   .o(edt_scan_out_buf_out[123]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_124_buf (.a(edt_scan_out[124]),
                                                                   .o(edt_scan_out_buf_out[124]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_125_buf (.a(edt_scan_out[125]),
                                                                   .o(edt_scan_out_buf_out[125]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_126_buf (.a(edt_scan_out[126]),
                                                                   .o(edt_scan_out_buf_out[126]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_127_buf (.a(edt_scan_out[127]),
                                                                   .o(edt_scan_out_buf_out[127]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_128_buf (.a(edt_scan_out[128]),
                                                                   .o(edt_scan_out_buf_out[128]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_129_buf (.a(edt_scan_out[129]),
                                                                   .o(edt_scan_out_buf_out[129]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_130_buf (.a(edt_scan_out[130]),
                                                                   .o(edt_scan_out_buf_out[130]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_131_buf (.a(edt_scan_out[131]),
                                                                   .o(edt_scan_out_buf_out[131]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_132_buf (.a(edt_scan_out[132]),
                                                                   .o(edt_scan_out_buf_out[132]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_133_buf (.a(edt_scan_out[133]),
                                                                   .o(edt_scan_out_buf_out[133]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_134_buf (.a(edt_scan_out[134]),
                                                                   .o(edt_scan_out_buf_out[134]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_135_buf (.a(edt_scan_out[135]),
                                                                   .o(edt_scan_out_buf_out[135]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_136_buf (.a(edt_scan_out[136]),
                                                                   .o(edt_scan_out_buf_out[136]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_137_buf (.a(edt_scan_out[137]),
                                                                   .o(edt_scan_out_buf_out[137]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_138_buf (.a(edt_scan_out[138]),
                                                                   .o(edt_scan_out_buf_out[138]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_139_buf (.a(edt_scan_out[139]),
                                                                   .o(edt_scan_out_buf_out[139]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_140_buf (.a(edt_scan_out[140]),
                                                                   .o(edt_scan_out_buf_out[140]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_141_buf (.a(edt_scan_out[141]),
                                                                   .o(edt_scan_out_buf_out[141]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_142_buf (.a(edt_scan_out[142]),
                                                                   .o(edt_scan_out_buf_out[142]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_143_buf (.a(edt_scan_out[143]),
                                                                   .o(edt_scan_out_buf_out[143]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_144_buf (.a(edt_scan_out[144]),
                                                                   .o(edt_scan_out_buf_out[144]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_145_buf (.a(edt_scan_out[145]),
                                                                   .o(edt_scan_out_buf_out[145]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_146_buf (.a(edt_scan_out[146]),
                                                                   .o(edt_scan_out_buf_out[146]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_147_buf (.a(edt_scan_out[147]),
                                                                   .o(edt_scan_out_buf_out[147]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_148_buf (.a(edt_scan_out[148]),
                                                                   .o(edt_scan_out_buf_out[148]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_149_buf (.a(edt_scan_out[149]),
                                                                   .o(edt_scan_out_buf_out[149]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_150_buf (.a(edt_scan_out[150]),
                                                                   .o(edt_scan_out_buf_out[150]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_151_buf (.a(edt_scan_out[151]),
                                                                   .o(edt_scan_out_buf_out[151]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_152_buf (.a(edt_scan_out[152]),
                                                                   .o(edt_scan_out_buf_out[152]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_153_buf (.a(edt_scan_out[153]),
                                                                   .o(edt_scan_out_buf_out[153]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_154_buf (.a(edt_scan_out[154]),
                                                                   .o(edt_scan_out_buf_out[154]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_155_buf (.a(edt_scan_out[155]),
                                                                   .o(edt_scan_out_buf_out[155]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_156_buf (.a(edt_scan_out[156]),
                                                                   .o(edt_scan_out_buf_out[156]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_157_buf (.a(edt_scan_out[157]),
                                                                   .o(edt_scan_out_buf_out[157]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_158_buf (.a(edt_scan_out[158]),
                                                                   .o(edt_scan_out_buf_out[158]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_159_buf (.a(edt_scan_out[159]),
                                                                   .o(edt_scan_out_buf_out[159]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_160_buf (.a(edt_scan_out[160]),
                                                                   .o(edt_scan_out_buf_out[160]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_161_buf (.a(edt_scan_out[161]),
                                                                   .o(edt_scan_out_buf_out[161]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_162_buf (.a(edt_scan_out[162]),
                                                                   .o(edt_scan_out_buf_out[162]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_163_buf (.a(edt_scan_out[163]),
                                                                   .o(edt_scan_out_buf_out[163]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_164_buf (.a(edt_scan_out[164]),
                                                                   .o(edt_scan_out_buf_out[164]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_165_buf (.a(edt_scan_out[165]),
                                                                   .o(edt_scan_out_buf_out[165]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_166_buf (.a(edt_scan_out[166]),
                                                                   .o(edt_scan_out_buf_out[166]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_167_buf (.a(edt_scan_out[167]),
                                                                   .o(edt_scan_out_buf_out[167]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_168_buf (.a(edt_scan_out[168]),
                                                                   .o(edt_scan_out_buf_out[168]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_169_buf (.a(edt_scan_out[169]),
                                                                   .o(edt_scan_out_buf_out[169]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_170_buf (.a(edt_scan_out[170]),
                                                                   .o(edt_scan_out_buf_out[170]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_171_buf (.a(edt_scan_out[171]),
                                                                   .o(edt_scan_out_buf_out[171]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_172_buf (.a(edt_scan_out[172]),
                                                                   .o(edt_scan_out_buf_out[172]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_173_buf (.a(edt_scan_out[173]),
                                                                   .o(edt_scan_out_buf_out[173]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_174_buf (.a(edt_scan_out[174]),
                                                                   .o(edt_scan_out_buf_out[174]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_175_buf (.a(edt_scan_out[175]),
                                                                   .o(edt_scan_out_buf_out[175]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_176_buf (.a(edt_scan_out[176]),
                                                                   .o(edt_scan_out_buf_out[176]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_177_buf (.a(edt_scan_out[177]),
                                                                   .o(edt_scan_out_buf_out[177]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_178_buf (.a(edt_scan_out[178]),
                                                                   .o(edt_scan_out_buf_out[178]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_179_buf (.a(edt_scan_out[179]),
                                                                   .o(edt_scan_out_buf_out[179]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_180_buf (.a(edt_scan_out[180]),
                                                                   .o(edt_scan_out_buf_out[180]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_181_buf (.a(edt_scan_out[181]),
                                                                   .o(edt_scan_out_buf_out[181]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_182_buf (.a(edt_scan_out[182]),
                                                                   .o(edt_scan_out_buf_out[182]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_183_buf (.a(edt_scan_out[183]),
                                                                   .o(edt_scan_out_buf_out[183]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_184_buf (.a(edt_scan_out[184]),
                                                                   .o(edt_scan_out_buf_out[184]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_185_buf (.a(edt_scan_out[185]),
                                                                   .o(edt_scan_out_buf_out[185]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_186_buf (.a(edt_scan_out[186]),
                                                                   .o(edt_scan_out_buf_out[186]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_187_buf (.a(edt_scan_out[187]),
                                                                   .o(edt_scan_out_buf_out[187]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_188_buf (.a(edt_scan_out[188]),
                                                                   .o(edt_scan_out_buf_out[188]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_189_buf (.a(edt_scan_out[189]),
                                                                   .o(edt_scan_out_buf_out[189]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_190_buf (.a(edt_scan_out[190]),
                                                                   .o(edt_scan_out_buf_out[190]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_191_buf (.a(edt_scan_out[191]),
                                                                   .o(edt_scan_out_buf_out[191]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_192_buf (.a(edt_scan_out[192]),
                                                                   .o(edt_scan_out_buf_out[192]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_193_buf (.a(edt_scan_out[193]),
                                                                   .o(edt_scan_out_buf_out[193]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_194_buf (.a(edt_scan_out[194]),
                                                                   .o(edt_scan_out_buf_out[194]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_195_buf (.a(edt_scan_out[195]),
                                                                   .o(edt_scan_out_buf_out[195]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_196_buf (.a(edt_scan_out[196]),
                                                                   .o(edt_scan_out_buf_out[196]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_197_buf (.a(edt_scan_out[197]),
                                                                   .o(edt_scan_out_buf_out[197]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_198_buf (.a(edt_scan_out[198]),
                                                                   .o(edt_scan_out_buf_out[198]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_199_buf (.a(edt_scan_out[199]),
                                                                   .o(edt_scan_out_buf_out[199]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_200_buf (.a(edt_scan_out[200]),
                                                                   .o(edt_scan_out_buf_out[200]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_201_buf (.a(edt_scan_out[201]),
                                                                   .o(edt_scan_out_buf_out[201]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_202_buf (.a(edt_scan_out[202]),
                                                                   .o(edt_scan_out_buf_out[202]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_203_buf (.a(edt_scan_out[203]),
                                                                   .o(edt_scan_out_buf_out[203]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_204_buf (.a(edt_scan_out[204]),
                                                                   .o(edt_scan_out_buf_out[204]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_205_buf (.a(edt_scan_out[205]),
                                                                   .o(edt_scan_out_buf_out[205]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_206_buf (.a(edt_scan_out[206]),
                                                                   .o(edt_scan_out_buf_out[206]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_207_buf (.a(edt_scan_out[207]),
                                                                   .o(edt_scan_out_buf_out[207]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_208_buf (.a(edt_scan_out[208]),
                                                                   .o(edt_scan_out_buf_out[208]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_209_buf (.a(edt_scan_out[209]),
                                                                   .o(edt_scan_out_buf_out[209]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_210_buf (.a(edt_scan_out[210]),
                                                                   .o(edt_scan_out_buf_out[210]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_211_buf (.a(edt_scan_out[211]),
                                                                   .o(edt_scan_out_buf_out[211]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_212_buf (.a(edt_scan_out[212]),
                                                                   .o(edt_scan_out_buf_out[212]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_213_buf (.a(edt_scan_out[213]),
                                                                   .o(edt_scan_out_buf_out[213]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_214_buf (.a(edt_scan_out[214]),
                                                                   .o(edt_scan_out_buf_out[214]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_215_buf (.a(edt_scan_out[215]),
                                                                   .o(edt_scan_out_buf_out[215]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_216_buf (.a(edt_scan_out[216]),
                                                                   .o(edt_scan_out_buf_out[216]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_217_buf (.a(edt_scan_out[217]),
                                                                   .o(edt_scan_out_buf_out[217]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_218_buf (.a(edt_scan_out[218]),
                                                                   .o(edt_scan_out_buf_out[218]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_219_buf (.a(edt_scan_out[219]),
                                                                   .o(edt_scan_out_buf_out[219]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_220_buf (.a(edt_scan_out[220]),
                                                                   .o(edt_scan_out_buf_out[220]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_221_buf (.a(edt_scan_out[221]),
                                                                   .o(edt_scan_out_buf_out[221]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_222_buf (.a(edt_scan_out[222]),
                                                                   .o(edt_scan_out_buf_out[222]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_223_buf (.a(edt_scan_out[223]),
                                                                   .o(edt_scan_out_buf_out[223]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_224_buf (.a(edt_scan_out[224]),
                                                                   .o(edt_scan_out_buf_out[224]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_225_buf (.a(edt_scan_out[225]),
                                                                   .o(edt_scan_out_buf_out[225]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_226_buf (.a(edt_scan_out[226]),
                                                                   .o(edt_scan_out_buf_out[226]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_227_buf (.a(edt_scan_out[227]),
                                                                   .o(edt_scan_out_buf_out[227]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_228_buf (.a(edt_scan_out[228]),
                                                                   .o(edt_scan_out_buf_out[228]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_229_buf (.a(edt_scan_out[229]),
                                                                   .o(edt_scan_out_buf_out[229]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_230_buf (.a(edt_scan_out[230]),
                                                                   .o(edt_scan_out_buf_out[230]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_231_buf (.a(edt_scan_out[231]),
                                                                   .o(edt_scan_out_buf_out[231]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_232_buf (.a(edt_scan_out[232]),
                                                                   .o(edt_scan_out_buf_out[232]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_233_buf (.a(edt_scan_out[233]),
                                                                   .o(edt_scan_out_buf_out[233]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_234_buf (.a(edt_scan_out[234]),
                                                                   .o(edt_scan_out_buf_out[234]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_235_buf (.a(edt_scan_out[235]),
                                                                   .o(edt_scan_out_buf_out[235]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_236_buf (.a(edt_scan_out[236]),
                                                                   .o(edt_scan_out_buf_out[236]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_237_buf (.a(edt_scan_out[237]),
                                                                   .o(edt_scan_out_buf_out[237]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_238_buf (.a(edt_scan_out[238]),
                                                                   .o(edt_scan_out_buf_out[238]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_239_buf (.a(edt_scan_out[239]),
                                                                   .o(edt_scan_out_buf_out[239]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_240_buf (.a(edt_scan_out[240]),
                                                                   .o(edt_scan_out_buf_out[240]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_241_buf (.a(edt_scan_out[241]),
                                                                   .o(edt_scan_out_buf_out[241]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_242_buf (.a(edt_scan_out[242]),
                                                                   .o(edt_scan_out_buf_out[242]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_243_buf (.a(edt_scan_out[243]),
                                                                   .o(edt_scan_out_buf_out[243]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_244_buf (.a(edt_scan_out[244]),
                                                                   .o(edt_scan_out_buf_out[244]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_245_buf (.a(edt_scan_out[245]),
                                                                   .o(edt_scan_out_buf_out[245]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_246_buf (.a(edt_scan_out[246]),
                                                                   .o(edt_scan_out_buf_out[246]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_247_buf (.a(edt_scan_out[247]),
                                                                   .o(edt_scan_out_buf_out[247]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_248_buf (.a(edt_scan_out[248]),
                                                                   .o(edt_scan_out_buf_out[248]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_249_buf (.a(edt_scan_out[249]),
                                                                   .o(edt_scan_out_buf_out[249]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_250_buf (.a(edt_scan_out[250]),
                                                                   .o(edt_scan_out_buf_out[250]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_251_buf (.a(edt_scan_out[251]),
                                                                   .o(edt_scan_out_buf_out[251]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_252_buf (.a(edt_scan_out[252]),
                                                                   .o(edt_scan_out_buf_out[252]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_253_buf (.a(edt_scan_out[253]),
                                                                   .o(edt_scan_out_buf_out[253]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_254_buf (.a(edt_scan_out[254]),
                                                                   .o(edt_scan_out_buf_out[254]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_255_buf (.a(edt_scan_out[255]),
                                                                   .o(edt_scan_out_buf_out[255]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_256_buf (.a(edt_scan_out[256]),
                                                                   .o(edt_scan_out_buf_out[256]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_257_buf (.a(edt_scan_out[257]),
                                                                   .o(edt_scan_out_buf_out[257]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_258_buf (.a(edt_scan_out[258]),
                                                                   .o(edt_scan_out_buf_out[258]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_259_buf (.a(edt_scan_out[259]),
                                                                   .o(edt_scan_out_buf_out[259]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_260_buf (.a(edt_scan_out[260]),
                                                                   .o(edt_scan_out_buf_out[260]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_261_buf (.a(edt_scan_out[261]),
                                                                   .o(edt_scan_out_buf_out[261]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_262_buf (.a(edt_scan_out[262]),
                                                                   .o(edt_scan_out_buf_out[262]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_263_buf (.a(edt_scan_out[263]),
                                                                   .o(edt_scan_out_buf_out[263]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_264_buf (.a(edt_scan_out[264]),
                                                                   .o(edt_scan_out_buf_out[264]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_265_buf (.a(edt_scan_out[265]),
                                                                   .o(edt_scan_out_buf_out[265]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_266_buf (.a(edt_scan_out[266]),
                                                                   .o(edt_scan_out_buf_out[266]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_267_buf (.a(edt_scan_out[267]),
                                                                   .o(edt_scan_out_buf_out[267]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_268_buf (.a(edt_scan_out[268]),
                                                                   .o(edt_scan_out_buf_out[268]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_269_buf (.a(edt_scan_out[269]),
                                                                   .o(edt_scan_out_buf_out[269]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_270_buf (.a(edt_scan_out[270]),
                                                                   .o(edt_scan_out_buf_out[270]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_271_buf (.a(edt_scan_out[271]),
                                                                   .o(edt_scan_out_buf_out[271]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_272_buf (.a(edt_scan_out[272]),
                                                                   .o(edt_scan_out_buf_out[272]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_273_buf (.a(edt_scan_out[273]),
                                                                   .o(edt_scan_out_buf_out[273]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_274_buf (.a(edt_scan_out[274]),
                                                                   .o(edt_scan_out_buf_out[274]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_275_buf (.a(edt_scan_out[275]),
                                                                   .o(edt_scan_out_buf_out[275]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_276_buf (.a(edt_scan_out[276]),
                                                                   .o(edt_scan_out_buf_out[276]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_277_buf (.a(edt_scan_out[277]),
                                                                   .o(edt_scan_out_buf_out[277]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_278_buf (.a(edt_scan_out[278]),
                                                                   .o(edt_scan_out_buf_out[278]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_279_buf (.a(edt_scan_out[279]),
                                                                   .o(edt_scan_out_buf_out[279]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_280_buf (.a(edt_scan_out[280]),
                                                                   .o(edt_scan_out_buf_out[280]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_281_buf (.a(edt_scan_out[281]),
                                                                   .o(edt_scan_out_buf_out[281]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_282_buf (.a(edt_scan_out[282]),
                                                                   .o(edt_scan_out_buf_out[282]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_283_buf (.a(edt_scan_out[283]),
                                                                   .o(edt_scan_out_buf_out[283]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_284_buf (.a(edt_scan_out[284]),
                                                                   .o(edt_scan_out_buf_out[284]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_285_buf (.a(edt_scan_out[285]),
                                                                   .o(edt_scan_out_buf_out[285]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_286_buf (.a(edt_scan_out[286]),
                                                                   .o(edt_scan_out_buf_out[286]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_287_buf (.a(edt_scan_out[287]),
                                                                   .o(edt_scan_out_buf_out[287]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_288_buf (.a(edt_scan_out[288]),
                                                                   .o(edt_scan_out_buf_out[288]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_289_buf (.a(edt_scan_out[289]),
                                                                   .o(edt_scan_out_buf_out[289]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_290_buf (.a(edt_scan_out[290]),
                                                                   .o(edt_scan_out_buf_out[290]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_291_buf (.a(edt_scan_out[291]),
                                                                   .o(edt_scan_out_buf_out[291]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_292_buf (.a(edt_scan_out[292]),
                                                                   .o(edt_scan_out_buf_out[292]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_293_buf (.a(edt_scan_out[293]),
                                                                   .o(edt_scan_out_buf_out[293]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_294_buf (.a(edt_scan_out[294]),
                                                                   .o(edt_scan_out_buf_out[294]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_295_buf (.a(edt_scan_out[295]),
                                                                   .o(edt_scan_out_buf_out[295]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_296_buf (.a(edt_scan_out[296]),
                                                                   .o(edt_scan_out_buf_out[296]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_297_buf (.a(edt_scan_out[297]),
                                                                   .o(edt_scan_out_buf_out[297]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_298_buf (.a(edt_scan_out[298]),
                                                                   .o(edt_scan_out_buf_out[298]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_299_buf (.a(edt_scan_out[299]),
                                                                   .o(edt_scan_out_buf_out[299]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_300_buf (.a(edt_scan_out[300]),
                                                                   .o(edt_scan_out_buf_out[300]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_301_buf (.a(edt_scan_out[301]),
                                                                   .o(edt_scan_out_buf_out[301]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_302_buf (.a(edt_scan_out[302]),
                                                                   .o(edt_scan_out_buf_out[302]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_303_buf (.a(edt_scan_out[303]),
                                                                   .o(edt_scan_out_buf_out[303]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_304_buf (.a(edt_scan_out[304]),
                                                                   .o(edt_scan_out_buf_out[304]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_305_buf (.a(edt_scan_out[305]),
                                                                   .o(edt_scan_out_buf_out[305]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_306_buf (.a(edt_scan_out[306]),
                                                                   .o(edt_scan_out_buf_out[306]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_307_buf (.a(edt_scan_out[307]),
                                                                   .o(edt_scan_out_buf_out[307]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_308_buf (.a(edt_scan_out[308]),
                                                                   .o(edt_scan_out_buf_out[308]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_309_buf (.a(edt_scan_out[309]),
                                                                   .o(edt_scan_out_buf_out[309]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_310_buf (.a(edt_scan_out[310]),
                                                                   .o(edt_scan_out_buf_out[310]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_311_buf (.a(edt_scan_out[311]),
                                                                   .o(edt_scan_out_buf_out[311]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_312_buf (.a(edt_scan_out[312]),
                                                                   .o(edt_scan_out_buf_out[312]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_313_buf (.a(edt_scan_out[313]),
                                                                   .o(edt_scan_out_buf_out[313]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_314_buf (.a(edt_scan_out[314]),
                                                                   .o(edt_scan_out_buf_out[314]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_315_buf (.a(edt_scan_out[315]),
                                                                   .o(edt_scan_out_buf_out[315]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_316_buf (.a(edt_scan_out[316]),
                                                                   .o(edt_scan_out_buf_out[316]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_317_buf (.a(edt_scan_out[317]),
                                                                   .o(edt_scan_out_buf_out[317]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_318_buf (.a(edt_scan_out[318]),
                                                                   .o(edt_scan_out_buf_out[318]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_319_buf (.a(edt_scan_out[319]),
                                                                   .o(edt_scan_out_buf_out[319]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_320_buf (.a(edt_scan_out[320]),
                                                                   .o(edt_scan_out_buf_out[320]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_321_buf (.a(edt_scan_out[321]),
                                                                   .o(edt_scan_out_buf_out[321]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_322_buf (.a(edt_scan_out[322]),
                                                                   .o(edt_scan_out_buf_out[322]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_323_buf (.a(edt_scan_out[323]),
                                                                   .o(edt_scan_out_buf_out[323]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_324_buf (.a(edt_scan_out[324]),
                                                                   .o(edt_scan_out_buf_out[324]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_325_buf (.a(edt_scan_out[325]),
                                                                   .o(edt_scan_out_buf_out[325]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_326_buf (.a(edt_scan_out[326]),
                                                                   .o(edt_scan_out_buf_out[326]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_327_buf (.a(edt_scan_out[327]),
                                                                   .o(edt_scan_out_buf_out[327]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_328_buf (.a(edt_scan_out[328]),
                                                                   .o(edt_scan_out_buf_out[328]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_329_buf (.a(edt_scan_out[329]),
                                                                   .o(edt_scan_out_buf_out[329]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_330_buf (.a(edt_scan_out[330]),
                                                                   .o(edt_scan_out_buf_out[330]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_331_buf (.a(edt_scan_out[331]),
                                                                   .o(edt_scan_out_buf_out[331]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_332_buf (.a(edt_scan_out[332]),
                                                                   .o(edt_scan_out_buf_out[332]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_333_buf (.a(edt_scan_out[333]),
                                                                   .o(edt_scan_out_buf_out[333]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_334_buf (.a(edt_scan_out[334]),
                                                                   .o(edt_scan_out_buf_out[334]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_335_buf (.a(edt_scan_out[335]),
                                                                   .o(edt_scan_out_buf_out[335]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_336_buf (.a(edt_scan_out[336]),
                                                                   .o(edt_scan_out_buf_out[336]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_337_buf (.a(edt_scan_out[337]),
                                                                   .o(edt_scan_out_buf_out[337]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_338_buf (.a(edt_scan_out[338]),
                                                                   .o(edt_scan_out_buf_out[338]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_339_buf (.a(edt_scan_out[339]),
                                                                   .o(edt_scan_out_buf_out[339]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_340_buf (.a(edt_scan_out[340]),
                                                                   .o(edt_scan_out_buf_out[340]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_341_buf (.a(edt_scan_out[341]),
                                                                   .o(edt_scan_out_buf_out[341]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_342_buf (.a(edt_scan_out[342]),
                                                                   .o(edt_scan_out_buf_out[342]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_343_buf (.a(edt_scan_out[343]),
                                                                   .o(edt_scan_out_buf_out[343]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_344_buf (.a(edt_scan_out[344]),
                                                                   .o(edt_scan_out_buf_out[344]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_345_buf (.a(edt_scan_out[345]),
                                                                   .o(edt_scan_out_buf_out[345]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_346_buf (.a(edt_scan_out[346]),
                                                                   .o(edt_scan_out_buf_out[346]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_347_buf (.a(edt_scan_out[347]),
                                                                   .o(edt_scan_out_buf_out[347]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_348_buf (.a(edt_scan_out[348]),
                                                                   .o(edt_scan_out_buf_out[348]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_349_buf (.a(edt_scan_out[349]),
                                                                   .o(edt_scan_out_buf_out[349]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_350_buf (.a(edt_scan_out[350]),
                                                                   .o(edt_scan_out_buf_out[350]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_351_buf (.a(edt_scan_out[351]),
                                                                   .o(edt_scan_out_buf_out[351]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_352_buf (.a(edt_scan_out[352]),
                                                                   .o(edt_scan_out_buf_out[352]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_353_buf (.a(edt_scan_out[353]),
                                                                   .o(edt_scan_out_buf_out[353]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_354_buf (.a(edt_scan_out[354]),
                                                                   .o(edt_scan_out_buf_out[354]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_355_buf (.a(edt_scan_out[355]),
                                                                   .o(edt_scan_out_buf_out[355]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_356_buf (.a(edt_scan_out[356]),
                                                                   .o(edt_scan_out_buf_out[356]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_357_buf (.a(edt_scan_out[357]),
                                                                   .o(edt_scan_out_buf_out[357]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_358_buf (.a(edt_scan_out[358]),
                                                                   .o(edt_scan_out_buf_out[358]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_359_buf (.a(edt_scan_out[359]),
                                                                   .o(edt_scan_out_buf_out[359]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_360_buf (.a(edt_scan_out[360]),
                                                                   .o(edt_scan_out_buf_out[360]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_361_buf (.a(edt_scan_out[361]),
                                                                   .o(edt_scan_out_buf_out[361]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_362_buf (.a(edt_scan_out[362]),
                                                                   .o(edt_scan_out_buf_out[362]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_363_buf (.a(edt_scan_out[363]),
                                                                   .o(edt_scan_out_buf_out[363]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_364_buf (.a(edt_scan_out[364]),
                                                                   .o(edt_scan_out_buf_out[364]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_365_buf (.a(edt_scan_out[365]),
                                                                   .o(edt_scan_out_buf_out[365]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_366_buf (.a(edt_scan_out[366]),
                                                                   .o(edt_scan_out_buf_out[366]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_367_buf (.a(edt_scan_out[367]),
                                                                   .o(edt_scan_out_buf_out[367]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_368_buf (.a(edt_scan_out[368]),
                                                                   .o(edt_scan_out_buf_out[368]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_369_buf (.a(edt_scan_out[369]),
                                                                   .o(edt_scan_out_buf_out[369]));
   i0sbfn000ab1n02x5 tessent_persistent_cell_edt_scan_out_370_buf (.a(edt_scan_out[370]),
                                                                   .o(edt_scan_out_buf_out[370]));

   firebird7_in_gate2_tessent_edt_intest_edt_decompressor firebird7_in_gate2_tessent_edt_intest_edt_decompressor_i (
      .edt_clock(edt_clock_buf_out),
      .edt_update(edt_update_buf_out),
      .edt_channels_in(edt_channels_out_from_controller),
      .edt_scan_in(edt_decompressor_out));

   firebird7_in_gate2_tessent_edt_intest_edt_compactor firebird7_in_gate2_tessent_edt_intest_edt_compactor_i (
      .edt_clock(edt_clock_buf_out),
      .edt_scan_out(edt_scan_out_buf_out),
      .masks_for_compactor_0(masks_for_compactor_0),
      .masks_for_compactor_1(masks_for_compactor_1),
      .edt_channels_out(edt_bypass_out));

   firebird7_in_gate2_tessent_edt_intest_edt_controller firebird7_in_gate2_tessent_edt_intest_edt_controller_i (
      .edt_clock(edt_clock_buf_out),
      .edt_update(edt_update_buf_out),
      .edt_low_power_shift_en(edt_low_power_shift_en_buf_out),
      .edt_channels_in(edt_channels_in_buf_out),
      .edt_decompressor_out(edt_decompressor_out),
      .edt_channels_out_from_controller(edt_channels_out_from_controller),
      .masks_for_compactor_0(masks_for_compactor_0),
      .masks_for_compactor_1(masks_for_compactor_1),
      .edt_scan_in(edt_bypass_in));

   firebird7_in_gate2_tessent_edt_intest_edt_bypass_logic firebird7_in_gate2_tessent_edt_intest_edt_bypass_logic_i (
      .edt_bypass(edt_bypass_buf_out),
      .edt_channels_in(edt_channels_in_buf_out),
      .edt_channels_out(edt_channels_out_buf_in),
      .edt_scan_in(edt_scan_in_buf_in),
      .edt_scan_out(edt_scan_out_buf_out),
      .edt_bypass_in(edt_bypass_in),
      .edt_bypass_out(edt_bypass_out));
endmodule


