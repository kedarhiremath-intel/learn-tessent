//
// Verilog format test patterns produced by Tessent Shell 2022.4
// Filename       : ./tsdb_outdir/patterns/firebird7_in_gate2.patterns_signoff/ICLNetwork.v
// Idstamp        : 2022.4:ec94:6099:0:0000
// Date           : Sun Nov  5 09:17:08 2023
//
// Begin_Verify_Section 
//   format            = Verilog 
//   top_module_name   = TB 
//   serial_flag       = OFF 
//   test_set_type     = IJTAG_TEST 
//   pad_value         = X 
//   one_setup         = ON 
//   no_initialization = ON 
// End_Verify_Section 
// Parameter File Keyword Settings 
//   SIM_CHANGE_PATH           true ; 
//   SIM_TOP_NAME              TB ; 
//   SIM_INSTANCE_NAME         DUT_inst ; 
//   SIM_CLOCK_MONITOR         true ; 
// End Parameter File Keyword Settings 


`define SIM_INSTANCE_NAME DUT_inst


`timescale 1ns / 100ps

module TB;

integer     _write_DIAG_file;
integer     _DIAG_file_header;
integer     _diag_file;
integer     _diag_chain_header;
integer     _diag_scan_header;
integer     _last_fail_pattern;
integer     _fail_pattern_cnt;
integer     _write_MASK_file;
integer     _MASK_file_header;
integer     _mask_file;
integer     _par_shift_cnt;
integer     _chain_test_;
integer     _compare_fail;
integer     _compare_fail_count;
integer     _compare_count;
integer     _compare_z_count;
integer     _bit_count;
integer     _report_bit_cnt;
integer     _miscompare_limit;
integer     _found_fail;
integer     _found_fail_per_cycle;
integer     _allow_bad_message_index;
integer     _end_vec_file_ok;
integer     _cycle_count, _save_cycle_count;
integer     _pattern_count, _repeat_count_nest[0:8], _repeat_count, _message_index;
integer     _index, _scan_index, _file_cnt, _max_index, _vec_pat_count, _save_index[0:8];
integer     _repeat_depth;
integer     _file_check;
integer     _run_testsetup;
integer     _in_testsetup;
integer     _start_pat;
integer     _end_pat;
integer     _end_after_setup;
integer     _no_setup;
integer     _save_state;
integer     _restart_state;
integer     _in_restart;
integer     _override_cfg;
integer     _in_range;
integer     _do_compare;
integer     _in_chaintest;
integer     _pat_num;
integer     _skipped_patterns;
integer     _end_simulation;
integer     _config_file;
integer     _fstat;
integer     _max_file_cnt;
reg[256*8:1] _vec_file_name;
reg[256*8:1] _cfg_file_name;
integer     _scan_shift_count;
reg[13:0]    _ibus;
reg[0:0]    _exp_obus, _msk_obus;
wire[0:0]   _sim_obus;
reg[2:0]    _pat_type;
reg         _tp_num;
reg         mgcdft_save_signal, mgcdft_restart_signal;
reg[38:0]   vect;

wire fdfx_powergood, secure_red, secure_orange, secure_insysbist, ijtag_tck, 
     ijtag_reset, ijtag_ce, ijtag_se, ijtag_ue, ijtag_sel, ijtag_si, 
     PD_TOP_bisr_shift_en, PD_TOP_bisr_clk, PD_TOP_bisr_reset, ijtag_so;

event       before_finish;
assign fdfx_powergood = _ibus[13];
assign secure_red = _ibus[12];
assign secure_orange = _ibus[11];
assign secure_insysbist = _ibus[10];
assign ijtag_tck = _ibus[9];
assign ijtag_reset = _ibus[8];
assign ijtag_ce = _ibus[7];
assign ijtag_se = _ibus[6];
assign ijtag_ue = _ibus[5];
assign ijtag_sel = _ibus[4];
assign ijtag_si = _ibus[3];
assign PD_TOP_bisr_shift_en = _ibus[2];
assign PD_TOP_bisr_clk = _ibus[1];
assign PD_TOP_bisr_reset = _ibus[0];

assign _sim_obus[0] = ijtag_so;

// Change Path Variables & Get Argument 
integer      _change_path; 
integer      _change_out_path; 
reg[512*8:1]  _new_path; 
reg[512*8:1]  _new_out_path; 
reg[512*8:1]  _new_filename; 
reg[512*8:1]  _vcd_dump_file_name; 
reg[512*8:1]  _utvcd_dump_file_name; 
reg[512*8:1]  _fsdb_dump_file_name; 
reg[512*8:1]  _qwave_dump_file_name; 
reg[512*8:1]  _tmp_filename; 
initial begin 
  _change_path = 0; 
  _change_out_path = 0; 
  if ($value$plusargs("NEWPATH=%s", _new_path)) begin 
    $display("Found New Path %0s\n", _new_path); 
    _change_path = 1; 
  end 
  if ($value$plusargs("NEWOUTPATH=%s", _new_out_path)) begin 
    $display("Found New Out Path %0s\n", _new_out_path); 
    _change_out_path = 1; 
  end 

`ifdef VCD
    $sformat(_vcd_dump_file_name, "ICLNetwork.v.dump");
    if(_change_out_path) begin 
      $sformat(_vcd_dump_file_name, "%0s/%0s", _new_out_path, _vcd_dump_file_name);
    end
    $dumpfile(_vcd_dump_file_name);
    $dumpvars;
`endif

`ifdef UTVCD
    $sformat(_utvcd_dump_file_name, "ICLNetwork.v.dump");
    if(_change_out_path) begin 
      $sformat(_utvcd_dump_file_name, "%0s/%0s", _new_out_path, _utvcd_dump_file_name);
    end
    $dumpfile(_utvcd_dump_file_name);
    $vtDump;
    $dumpvars;
`endif

`ifdef debussy
    $sformat(_fsdb_dump_file_name, "ICLNetwork.v.fsdb");
    if(_change_out_path) begin 
      $sformat(_fsdb_dump_file_name, "%0s/%0s", _new_out_path, _fsdb_dump_file_name);
    end
    $fsdbDumpfile(_fsdb_dump_file_name);
    $fsdbDumpvars;
`endif

`ifdef QWAVE
    $sformat(_qwave_dump_file_name, "ICLNetwork.v.qwave.db");
    if(_change_out_path) begin 
      $sformat(_qwave_dump_file_name, "%0s/%0s", _new_out_path, _qwave_dump_file_name);
    end
    $qwavedb_dumpvars_filename(_qwave_dump_file_name);
    $qwavedb_dumpvars;
`endif
end 

reg /* sparse */[63:0] _nam_obus[0:0];
initial begin 
   if(_change_path) begin 
     $sformat(_new_filename,"%0s/ICLNetwork.v.po.name",_new_path); 
     $display("Loading %0s\n", _new_filename ); 
     $readmemh(_new_filename,_nam_obus,0,0); 
   end 
   else begin
     $display("Loading ICLNetwork.v.po.name");
     $readmemh("ICLNetwork.v.po.name",_nam_obus,0,0);
   end 
end 


// Declare Wires for tracking Vector Type
reg[3:0] _MGCDFT_VECTYPE ;
reg[160:0] _procedure_string ;
reg mgcdft_test_setup, mgcdft_load_unload, mgcdft_shift,
     mgcdft_single_shift, mgcdft_shift_extra, 
     mgcdft_shadow_control, mgcdft_master_observe,
     mgcdft_shadow_observe, mgcdft_skew_load, 
     mgcdft_seq_transparent, mgcdft_launch_capture,
     mgcdft_clock_proc, mgcdft_test_end, mgcdft_unknown; 

event       set_vector_type;
always @(_MGCDFT_VECTYPE) begin
  assign mgcdft_test_setup      = 1'b0;
  assign mgcdft_load_unload     = 1'b0;
  assign mgcdft_shift           = 1'b0;
  assign mgcdft_single_shift    = 1'b0;
  assign mgcdft_shift_extra     = 1'b0;
  assign mgcdft_shadow_control  = 1'b0;
  assign mgcdft_master_observe  = 1'b0;
  assign mgcdft_shadow_observe  = 1'b0;
  assign mgcdft_skew_load       = 1'b0;
  assign mgcdft_seq_transparent = 1'b0;
  assign mgcdft_launch_capture  = 1'b0;
  assign mgcdft_clock_proc      = 1'b0;
  assign mgcdft_test_end        = 1'b0;
  assign mgcdft_unknown         = 1'b0;
  case (_MGCDFT_VECTYPE)
    4'b0001: begin
               assign mgcdft_test_setup      = 1'b1;
               _procedure_string = "TEST_SETUP";
               _scan_shift_count = 0;
             end
    4'b0010: begin
               assign mgcdft_load_unload     = 1'b1;
               _procedure_string = "LOAD";
               _scan_shift_count = 0;
             end
    4'b0011: begin
               assign mgcdft_shift           = 1'b1;
               _procedure_string = "SHIFT";
               if(!(_scan_shift_count)) begin
                 _scan_shift_count = 1;
               end
             end
    4'b0100: begin
               assign mgcdft_single_shift    = 1'b1;
               _procedure_string = "SINGLE_SHIFT";
               if(!(_scan_shift_count)) begin
                 _scan_shift_count = 1;
               end
             end
    4'b0101: begin
               assign mgcdft_shift_extra     = 1'b1;
               _procedure_string = "SHIFT_EXTRA";
               _scan_shift_count = 0;
             end
    4'b0110: begin
               assign mgcdft_shadow_control  = 1'b1;
               _procedure_string = "SHADOW_CONTROL";
               _scan_shift_count = 0;
             end
    4'b0111: begin
               assign mgcdft_master_observe  = 1'b1;
               _procedure_string = "MASTER_OBSERVE";
               _scan_shift_count = 0;
             end
    4'b1000: begin
               assign mgcdft_shadow_observe  = 1'b1;
               _procedure_string = "SHADOW_OBSERVE";
               _scan_shift_count = 0;
             end
    4'b1001: begin
               assign mgcdft_skew_load       = 1'b1;
               _procedure_string = "SKEW_LOAD";
               _scan_shift_count = 0;
             end
    4'b1010: begin
               assign mgcdft_seq_transparent = 1'b1;
               _procedure_string = "SEQ_TRANSPARENT";
               _scan_shift_count = 0;
             end
    4'b1011: begin
               assign mgcdft_launch_capture  = 1'b1;
               _procedure_string = "LAUNCH_CAPTURE";
               _scan_shift_count = 0;
             end
    4'b1101: begin
               assign mgcdft_clock_proc      = 1'b1;
               _procedure_string = "CLOCK_PROC";
               _scan_shift_count = 0;
             end
    4'b1111: begin
               assign mgcdft_test_end        = 1'b1;
               _procedure_string = "TEST_END";
               _scan_shift_count = 0;
             end
    4'b0000: begin
               assign mgcdft_unknown         = 1'b1;
               _procedure_string = "UNKNOWN";
               _scan_shift_count = 0;
             end
    default: begin
               assign mgcdft_unknown         = 1'b1;
               _procedure_string = "UNKNOWN";
               _scan_shift_count = 0;
             end
  endcase
end

function integer do_finish_summary;
input local_end_vec_file_ok;
integer local_end_vec_file_ok;
begin
  if (_end_vec_file_ok) begin
     $display("\nSimulation finished at time %.0f", $realtime);
     $display("Number of miscompares            = %d", _compare_fail_count);
     $display("Number of 0/1 compares           = %d", _compare_count);
     $display("Number of Z compares             = %d\n", _compare_z_count);
  end

  if ((_end_vec_file_ok) && (_compare_fail == 0) && (_compare_fail_count == 0)) begin
     $display("No error between simulated and expected patterns\n");
  end

  if ((_compare_fail != 0) || (_compare_fail_count != 0)) begin
     $display("Error between simulated and expected patterns\n");
  end

do_finish_summary = local_end_vec_file_ok;
end
endfunction


event       compare_exp_sim_obus;
always @(compare_exp_sim_obus) begin
 _found_fail = 0;
 if (_do_compare) begin
 for(_bit_count = 0;
     (_bit_count < 1);
      _bit_count =_bit_count +1) begin
   if (_msk_obus[_bit_count] === 1'b1) begin
     if (_exp_obus[_bit_count] === 1'bZ) begin
       _compare_z_count = _compare_z_count + 1;
     end
     else begin
       _compare_count = _compare_count + 1;
     end
   end
 end
  if (_exp_obus !== _sim_obus) begin
     for(_bit_count = 0;
         ((_bit_count < 1)&&(_found_fail==0));
          _bit_count =_bit_count +1) begin
        if ((_msk_obus[_bit_count] === 1'b1) &&
            (_exp_obus[_bit_count] !== _sim_obus[_bit_count])) begin
           _found_fail = 1;
           _found_fail_per_cycle = 1;
        end
     end
  end
  if (_found_fail == 1) begin
     for(_bit_count = 0;
         ((_bit_count < 1)&&((_miscompare_limit==0)||(_compare_fail<=_miscompare_limit)));
          _bit_count =_bit_count +1) begin
      if ((_msk_obus[_bit_count] === 1'b1) &&
          (_exp_obus[_bit_count] !== _sim_obus[_bit_count])) begin
        _compare_fail_count = _compare_fail_count + 1;
        $write($realtime, "ns: Mismatch at pin %d name %s, Simulated %b, Expected %b\n",_bit_count,_nam_obus[_bit_count],_sim_obus[_bit_count],_exp_obus[_bit_count]);
        if (_write_DIAG_file == 1) begin
          if (_DIAG_file_header == 0) begin
            if ((_start_pat > -1) && (_end_pat > -1)) begin
              $sformat(_tmp_filename, "ICLNetwork.v_%0d_%0d.fail",
                       _start_pat, _end_pat);
            end
            else if (_start_pat > -1) begin
              $sformat(_tmp_filename, "ICLNetwork.v_%0d.fail",
                       _start_pat);
            end
            else if (_end_pat > -1) begin
              $sformat(_tmp_filename, "ICLNetwork.v__%0d.fail",
                       _end_pat);
            end
            else begin
              $sformat(_tmp_filename, "ICLNetwork.v.fail");
            end
            if(_change_out_path) begin 
              $sformat(_tmp_filename, "%0s/%0s", _new_out_path, _tmp_filename);
            end
            _diag_file = $fopen(_tmp_filename);
            if (_diag_file == 0) begin
              $display("ERROR: Couldn't open .fail file %0s, simulation aborted\n", _tmp_filename);
              ->before_finish;
              #0;
              $finish;
            end
            if(_change_out_path) begin 
              $fwrite(_diag_file, "// This File is simulation generated (%0s/ICLNetwork.v)\n", _new_out_path);
            end
            else begin
              $fwrite(_diag_file, "// This File is simulation generated (ICLNetwork.v)\n");
            end
            $fwrite(_diag_file, "format cycle\n");
            $fwrite(_diag_file, " failures_begin\n");
            $fwrite(_diag_file, "//cycle_number  PO_name  expected_value  simulated_value  ");
            $fwrite(_diag_file, "pattern_id  chain_name  cell_number\n\n");
            _DIAG_file_header = 1;
          end
          if ((_pattern_count == _last_fail_pattern) && (_pattern_count == 0)) begin
             _fail_pattern_cnt = 1; 
          end
          if (_pattern_count > _last_fail_pattern) begin 
             _fail_pattern_cnt = _fail_pattern_cnt + 1;
             _last_fail_pattern = _pattern_count;
          end

          $fwrite(_diag_file, "%d  %s ", _cycle_count, _nam_obus[_bit_count]);
          case ( _exp_obus[_bit_count] )
            1'b1: begin
                    $fwrite(_diag_file, "            H"); 
                  end
            1'b0: begin
                    $fwrite(_diag_file, "            L"); 
                  end
            1'bZ: begin
                    $fwrite(_diag_file, "            Z"); 
                  end
          endcase
          case ( _sim_obus[_bit_count] )
            1'b1: begin
                    $fwrite(_diag_file, " H  // Pattern %d ", _pattern_count); 
                  end
            1'b0: begin
                    $fwrite(_diag_file, " L  // Pattern %d ", _pattern_count); 
                  end
            1'bZ: begin
                    $fwrite(_diag_file, " Z  // Pattern %d ", _pattern_count); 
                  end
            1'bX: begin
                    $fwrite(_diag_file, " X  // Pattern %d ", _pattern_count); 
                  end
          endcase
         if (_scan_shift_count == 0) begin
                 $fwrite(_diag_file, ", simulation_time=%.0f\n", $realtime);
         end // EndIf  _ScanShift_count
        end // EndIf _write_DIAG_file
        if (_write_MASK_file == 1) begin
          if (_MASK_file_header == 0) begin
            if ((_start_pat > -1) && (_end_pat > -1)) begin
              $sformat(_tmp_filename, "ICLNetwork.v_%0d_%0d.mask",
                       _start_pat, _end_pat);
            end
            else if (_start_pat > -1) begin
              $sformat(_tmp_filename, "ICLNetwork.v_%0d.mask",
                       _start_pat);
            end
            else if (_end_pat > -1) begin
              $sformat(_tmp_filename, "ICLNetwork.v__%0d.mask",
                       _end_pat);
            end
            else begin
              $sformat(_tmp_filename, "ICLNetwork.v.mask");
            end
            if(_change_out_path) begin 
              $sformat(_tmp_filename, "%0s/%0s", _new_out_path, _tmp_filename);
            end
            _mask_file = $fopen(_tmp_filename);
            if (_mask_file == 0) begin
              $display("ERROR: Couldn't open .mask file %0s, simulation aborted\n", _tmp_filename);
              ->before_finish;
              #0;
              $finish;
            end
            $fwrite(_mask_file, "%s\n%s\n", "type mask", "");
            _MASK_file_header = 1;
          end
          if (_chain_test_ == 0) begin
            $fwrite(_mask_file, "%d %s\n", _pattern_count,_nam_obus[_bit_count]);
          end
          if (_chain_test_ == 1) begin
            $fwrite(_mask_file, "// %d %s\n", _pattern_count,_nam_obus[_bit_count]);
          end
        end
      end
    end
    _compare_fail = _compare_fail + 1;
  end
 end // if _do_compare
end

reg[38:0]     mem [0:3441479];
firebird7_in DUT_inst (.fdfx_powergood(fdfx_powergood), 
     .secure_red(secure_red), .secure_orange(secure_orange), 
     .secure_insysbist(secure_insysbist), .ijtag_tck(ijtag_tck), 
     .ijtag_reset(ijtag_reset), .ijtag_ce(ijtag_ce), 
     .ijtag_se(ijtag_se), .ijtag_ue(ijtag_ue), 
     .ijtag_sel(ijtag_sel), .ijtag_si(ijtag_si), 
     .PD_TOP_bisr_shift_en(PD_TOP_bisr_shift_en), 
     .PD_TOP_bisr_clk(PD_TOP_bisr_clk), 
     .PD_TOP_bisr_reset(PD_TOP_bisr_reset), .ijtag_so(ijtag_so));

initial begin
_in_restart = 0;
while (_in_restart < 2) begin
_in_restart = _in_restart + 1;
_restart_state     = -1;
if ($value$plusargs("RESTART=%d", _restart_state)) begin
  $display(" Found RESTART   %d", _restart_state);
end

if ((_in_restart < 2) || (_restart_state == 1)) begin
mgcdft_save_signal = 1'b0;
mgcdft_restart_signal = 1'b0;
if (_restart_state == 1) begin
  #0;
  mgcdft_restart_signal = 1'b1;
//  $display("Reading checkpoint ICLNetwork.v.dat");
//  $restart("ICLNetwork.v.dat");
end

#0;
mgcdft_save_signal = 1'b0;
mgcdft_restart_signal = 1'b0;
_compare_fail = 0;
_compare_fail_count = 0;
_compare_count = 0;
_compare_z_count = 0;
_pattern_count = 0;
_cycle_count = 0;
_save_cycle_count = 0;
_write_DIAG_file = 0; // change to 1, to generate file
_write_MASK_file = 0; // change to 1, to generate file
_DIAG_file_header = 0;
_diag_file = 0;
_diag_chain_header = 0;
_diag_scan_header = 0;
_fail_pattern_cnt = 0;
_last_fail_pattern = 0;
_MASK_file_header = 0;
_mask_file = 0;
_chain_test_ = 0;
_par_shift_cnt = 0;
_report_bit_cnt = 0;
// Limit # of miscompares before aborting simulation (non-zero)
_miscompare_limit = 0; 
_end_vec_file_ok = 0; 
_scan_shift_count = 0;
_run_testsetup  = 0;
_in_testsetup = 0;
_start_pat      = -1;
_end_pat        = -1;
_end_after_setup = -1;
_no_setup       = -1;
_save_state     = -1;
_override_cfg   = 0;
_pat_num        = -1;
_in_range       = 1;
_do_compare     = 1;
_in_chaintest   = 0;

_skipped_patterns = 0;

_end_simulation   = 0;

if ($value$plusargs("STARTPAT=%d", _start_pat)) begin
  if (_start_pat > -1) begin
    $display(" Found Start pattern number %d", _start_pat);
    _in_range = 0;
    _do_compare = 0;
  end
  else begin
    $display(" Ignoring negative Start pattern number   %d", _start_pat);
    _start_pat = -1;
  end
end
if ($value$plusargs("ENDPAT=%d", _end_pat)) begin
  if (_end_pat > -1) begin
    $display(" Found End pattern number   %d", _end_pat);
  end
  else begin
    $display(" Ignoring negative End pattern number   %d", _end_pat);
    _end_pat = -1;
  end
end

if ($value$plusargs("CHAINTEST=%d", _in_chaintest)) begin
  if (_in_chaintest) begin
    $display(" Found ChainTest identifier %d", _in_chaintest);
  end
end

if ($value$plusargs("END_AFTER_SETUP=%d", _end_after_setup)) begin
  $display(" Found End after setup   %d", _end_after_setup);
  if (_end_after_setup > 0) begin
    _end_pat = 0;
    _in_chaintest = 1;
  end
end

if ($value$plusargs("SKIP_SETUP=%d", _no_setup)) begin
  $display(" Found Skip setup   %d", _no_setup);
  if (_no_setup > 0) begin
    if (_start_pat == -1) begin
      _start_pat = 0;
      _in_chaintest = 1;
    end
    _run_testsetup = 0;
    _in_range = 0;
    _do_compare = 0;
  end
end

if ($value$plusargs("SAVE=%d", _save_state)) begin
  $display(" Found SAVE   %d", _save_state);
end

if ($value$plusargs("CONFIG=%0s", _cfg_file_name)) begin
  $display(" Found CONFIG identifier   %0s", _cfg_file_name);
  _override_cfg = 1;
end
else begin
  _cfg_file_name = "ICLNetwork.v.cfg";
end

if ((_end_pat != -1) && (_end_pat < _start_pat)) begin
  _start_pat = -1;
  _in_range = 1;
  _do_compare = 1;
  $display("STARTPAT less than ENDPAT, ignoring STARTPAT ");
end
_allow_bad_message_index = 0;
if ($value$plusargs("ALLOW_BAD_MESSAGE_INDEX=%d", _allow_bad_message_index)) begin
  $display(" Found ALLOW_BAD_MESSAGE_INDEX %d", _allow_bad_message_index);
end

// read vector config file
if(_override_cfg) begin 
  _config_file = $fopen(_cfg_file_name, "r");
end
else begin
if(_change_path) begin 
  $sformat(_new_filename,"%0s/ICLNetwork.v.cfg",_new_path); 
  _config_file = $fopen(_new_filename, "r");
end
else begin
  _config_file = $fopen("ICLNetwork.v.cfg", "r");
end

end

if (_config_file == 0) begin
  $display("ERROR: Couldn't open configuration file, simulation aborted\n");
  ->before_finish;
  #0;
  $finish;
end
_fstat = 0;
if (_start_pat != -1) begin
  if (_no_setup > 0) begin
  $display("BEGIN pattern read loop  Skip test_setup\n");
  end
  else if (_in_chaintest == 0) begin
    if (_end_pat != -1) begin
    $display("BEGIN pattern read loop  Start pattern (%d) End pattern (%d)\n",
_start_pat,_end_pat);
    end
    else begin
    $display("BEGIN pattern read loop  Start pattern (%d) \n",
_start_pat);
    end
  end
  else begin
    if (_end_pat != -1) begin
    $display("BEGIN pattern read loop  Start chain pattern (%d) End chain pattern (%d)\n",
_start_pat,_end_pat);
    end
    else begin
    $display("BEGIN pattern read loop  Start chain pattern (%d)\n",
_start_pat);
    end
  end
end
else if (_end_pat != -1) begin
  if (_end_after_setup > 0) begin
  $display("BEGIN pattern read loop  End after test_setup\n");
  end
  else if (_in_chaintest == 0) begin
  $display("BEGIN pattern read loop  End pattern (%d)\n", _end_pat);
  end
  else begin
  $display("BEGIN pattern read loop  End chain pattern (%d)\n", _end_pat);
  end
end

// begin pattern read loop
while (!$feof(_config_file) && (!_end_simulation))
begin
         _fstat = $fscanf(_config_file, "%s", _vec_file_name);
         _fstat = $fscanf(_config_file, "%d", _max_index);
   if (_fstat != -1) begin
         _fstat = $fscanf(_config_file, "%d", _vec_pat_count);
         if (_fstat == -1) begin
           _vec_pat_count = -1;
         end
         // skip .vec file if _start_pat greater than this
         if ((_start_pat != -1) && !_in_range && (_vec_pat_count != -1) &&
             !_in_testsetup && !_in_chaintest &&
             ((_pat_num + _vec_pat_count) < _start_pat)) begin
           _max_index = -1;
           if (_chain_test_) begin
             _pattern_count = 0;
             _pat_num = 0;
           end
           _pat_num = _pat_num + _vec_pat_count;
           _skipped_patterns = _skipped_patterns + _vec_pat_count;
           _end_vec_file_ok = 1;
           _chain_test_ = 0;
            $display("Skipping %0s\n", _vec_file_name);
         end
         else begin
          if(_change_path) begin 
            $sformat(_new_filename,"%0s/%0s",_new_path, _vec_file_name); 
            $display("Loading %0s\n", _new_filename ); 
            $readmemb(_new_filename, mem, 0, _max_index);
         end
         else begin
           $display("Loading %0s\n", _vec_file_name);
           $readmemb(_vec_file_name, mem, 0, _max_index);
         end
           _end_vec_file_ok = 0;
         end
   end
   else begin
     _max_index = -1;
     _vec_pat_count = -1;
   end
   _scan_index = 0;
   _repeat_count_nest[0] = 0;
   _repeat_count = 0;
   _repeat_depth = 0;
   _message_index = 0;
   _save_index[0] = 0;
   for (_index=0; _index <= _max_index; _index = _index+1)
   begin
      vect = mem[_index];
      _exp_obus=1'bX;
      _msk_obus=1'b0;
      _MGCDFT_VECTYPE = vect[3:0];
      _pat_type = vect[6:4];
      _tp_num = vect[7];
      //    Range Check
      if ((_start_pat != -1) && ((_start_pat != 0) || (!_in_testsetup)) &&
          ((!_chain_test_)||(_chain_test_ && _in_chaintest))) begin
        if (!_chain_test_ && _in_chaintest && !_in_range && !_in_testsetup) begin
          _in_range = 1;
          _do_compare = 1;
        end
        if ((_pat_num == _start_pat) && !_in_range) begin
          _in_range = 1;
          _do_compare = 0;
          _pattern_count = (_pat_num - 1);
          if (_pattern_count < 0) begin
            _pattern_count = 0;
          end
        end
        if (_pat_num == (_start_pat + 1)) begin
          _do_compare = 1;
        end
      end

      if ((_end_pat != -1) && (_pattern_count > _end_pat) && 
          ((!_chain_test_)||(_chain_test_ && _in_chaintest))) begin
         // simulation complete, exit
         _index = _max_index + 1;
         _end_vec_file_ok = 1;
         _end_simulation = 1;
      end
      if ((_index > 0) && (_end_pat != -1) && !_chain_test_ && _in_chaintest &&
          !_run_testsetup) begin
         // simulation complete, exit
         _index = _max_index + 1;
         _end_vec_file_ok = 1;
         _end_simulation = 1;
      end
      if ((_in_range) || (_run_testsetup)) begin
      case (_pat_type)
         3'b000:  begin // end vector
            _index = _max_index + 1;
         end // end vector
         3'b001: ;// skip scan vector, handled by shift vector
         3'b010:  begin // broadside vector
            _found_fail_per_cycle = 0;
            if (vect[8] == 1'b1) begin
               _pattern_count = _pattern_count + 1;
               _par_shift_cnt = 0;
              if ((!_do_compare) && (_pattern_count >= _start_pat)) begin
                _do_compare = 1;
              end
              if ((_end_pat != -1) && (_pattern_count > _end_pat) && 
                  ((!_chain_test_)||(_chain_test_ && _in_chaintest))) begin
                // simulation complete, exit
                _index = _max_index + 1;
                _end_vec_file_ok = 1;
                _end_simulation = 1;
                _in_range = 0;
              end
            end
            if (vect[8] === 1'bz) begin
               _pattern_count = 0;
               _par_shift_cnt = 0;
            end
            if(_scan_shift_count) begin
               _scan_shift_count = _scan_shift_count + 1;
            end
            case (_tp_num)
               1'b1: begin // timeplate 1 - gen_tp1
                  _ibus[9] = 1'b0;
                  _ibus[1] = 1'b0;
                  _ibus[13:10] = vect[24:21];
                  _ibus[8] = vect[19];
                  _ibus[3] = vect[14];
                  _ibus[0] = vect[11];

                  #24; // 24 ns
                  _exp_obus[0] = vect[10];
                  _msk_obus[0] = vect[9];
                  #0;
                  ->compare_exp_sim_obus;
                  if ((_miscompare_limit)&&(_compare_fail>=_miscompare_limit)) begin
                    $display("ERROR: exceeded miscompare limit(%d), exiting simulation",_miscompare_limit);
                    _end_vec_file_ok = 1;
                    if (_DIAG_file_header == 1) begin
                       if (_diag_scan_header==1) begin
                         $fwrite(_diag_file, "last_pattern_applied %d\n", _pattern_count);
                       end
                       $fwrite(_diag_file, "// failing_patterns=%d simulated_patterns=%d", _fail_pattern_cnt, (_pattern_count+1));
                       $fwrite(_diag_file, " simulation_time=", $realtime, ";\n");
                       $fwrite(_diag_file, "failure_file_end\n");
                       $fclose(_diag_file);
                    end
                    _end_vec_file_ok = do_finish_summary(_end_vec_file_ok);
                    ->before_finish;
                    #0;
                    $finish;
                  end

                  #1; // 25 ns
                  _ibus[9] = vect[20];
                  _ibus[1] = vect[12];

                  #24; // 49 ns
                  _ibus[5] = vect[16];

                  #26; // 75 ns
                  _ibus[9] = 1'b0;
                  _ibus[1] = 1'b0;

                  #24; // 99 ns
                  _ibus[7:6] = vect[18:17];
                  _ibus[4] = vect[15];
                  _ibus[2] = vect[13];

                  #1; // 100 ns
               end // timeplate 1 - gen_tp1
               default: begin
                  $display("ERROR: corrupt timeplate number\n");
                  ->before_finish;
                  #0;
                  $finish;
               end
            endcase // _tp_num
            _cycle_count = _cycle_count + 1;
            _par_shift_cnt = 0;
         end // broadside vector
         3'b011:  begin // status message vector
            _message_index = vect[38:7];
            case (_message_index)
               0: begin
                  $display("Begin chain test\n");
                 _chain_test_ = 1;
                  _diag_chain_header = 0;
               end
               1: begin
                 _chain_test_ = 0;
                  if (_diag_chain_header) begin
                    $fwrite(_diag_file, "last_pattern_applied %d\n", _pattern_count);
                  end
                  _diag_scan_header = 0;
                  if ((_start_pat > -1) || (_end_pat > -1)) begin
                    if (_pat_num > -1) begin
                        $display("Simulated chain pattern %d\n",_pat_num);
                    end
                  end
                  _pat_num = -1;
                  _pattern_count = 0;
                  $display("End chain test\n");
               end
               2: begin
                  $display("Status update: simulated through pattern %d\n",_pattern_count);
               end
               3: begin
                  _end_vec_file_ok = 1;
                  if ((_start_pat > -1) || (_end_pat > -1)) begin
                    if (_pat_num > -1) begin
                      if (!_chain_test_) begin
                        $display("Simulated pattern %d\n",_pat_num);
                      end
                    end
                  end
               end
               4: begin // start of atpg pattern
                  if ((_start_pat > -1) || (_end_pat > -1)) begin
                    if (_pat_num > -1) begin
                      if (_chain_test_) begin
                        $display("Simulated chain pattern %d\n",_pat_num);
                      end
                      else begin
                        $display("Simulated pattern %d\n",_pat_num);
                      end
                    end
                  end
                  _pat_num = _pat_num + 1;
                  _run_testsetup  = 0;
                  _in_testsetup  = 0;
                  if (_end_after_setup  > 0) begin
                    //simulation complete, exit
                    _index = _max_index + 1;
                    _end_vec_file_ok = 1;
                    _end_simulation = 1;
                    _in_range = 0;
                  end
               end
               20: begin
                  $display($realtime, "ns: Pattern_set firebird7_in");
               end
               21: begin
                  $display($realtime, "ns:  Activate selection of the following scan muxes:");
               end
               22: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               23: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               24: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               25: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.scan_in_mux, selection 1: sib, ltest_en = 2'bxx -> scan_in_mux = ijtag_si");
               end
               26: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               27: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               28: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               29: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               30: begin
                  $display($realtime, "ns:  Scan in verification pattern to the following scan registers:");
               end
               31: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.sib, load value = 1");
               end
               32: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.sib, load value = 1");
               end
               33: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.sib, load value = 0");
               end
               34: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.sib, load value = 0");
               end
               35: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.sib, load value = 1");
               end
               36: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.sib, load value = 1");
               end
               37: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.sib, load value = 0");
               end
               38: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_inst.sib, load value = 1");
               end
               39: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_sri_inst.sib ");
                  end
               end
               40: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.sib ");
                  end
               end
               41: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.sib ");
                  end
               end
               42: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_sti_inst.sib ");
                  end
               end
               43: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_spare_inst.sib ");
                  end
               end
               44: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_upm_inst.sib ");
                  end
               end
               45: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.sib ");
                  end
               end
               46: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.sib ");
                  end
               end
               47: begin
                  $display($realtime, "ns:  Scan out verification pattern from the following scan registers:");
               end
               48: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.sib, expected value = 1");
               end
               49: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.sib, expected value = 1");
               end
               50: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.sib, expected value = 0");
               end
               51: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.sib, expected value = 0");
               end
               52: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.sib, expected value = 1");
               end
               53: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.sib, expected value = 1");
               end
               54: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.sib, expected value = 0");
               end
               55: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_inst.sib, expected value = 1");
               end
               56: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               57: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_sri_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               58: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_sri_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               59: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_local_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               60: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_ctrl_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               61: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_edt_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               62: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               63: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               64: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.sib, load value = 0");
               end
               65: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.sib, load value = 0");
               end
               66: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.sib, load value = 1");
               end
               67: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.sib, load value = 1");
               end
               68: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.sib, load value = 0");
               end
               69: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.sib, load value = 0");
               end
               70: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_edt_inst.sib, load value = 1");
               end
               71: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_ctrl_inst.sib, load value = 1");
               end
               72: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_local_inst.sib, load value = 0");
               end
               73: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_sri_local_inst.sib ");
                  end
               end
               74: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_sri_ctrl_inst.sib ");
                  end
               end
               75: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_edt_inst.sib ");
                  end
               end
               76: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_occ_inst.sib ");
                  end
               end
               77: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_sib_ssn_inst.sib ");
                  end
               end
               78: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.sib, expected value = 0");
               end
               79: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.sib, expected value = 0");
               end
               80: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.sib, expected value = 1");
               end
               81: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.sib, expected value = 1");
               end
               82: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.sib, expected value = 0");
               end
               83: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.sib, expected value = 0");
               end
               84: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_edt_inst.sib, expected value = 1");
               end
               85: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_ctrl_inst.sib, expected value = 1");
               end
               86: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_local_inst.sib, expected value = 0");
               end
               87: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_local_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               88: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.sib, load value = 1");
               end
               89: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.sib, load value = 0");
               end
               90: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.sib, load value = 0");
               end
               91: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.sib, load value = 1");
               end
               92: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.sib, load value = 1");
               end
               93: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr4_inst.tdr[0:0], load value = 0");
               end
               94: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr3_inst.tdr[0:0], load value = 0");
               end
               95: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr2_inst.tdr[0:0], load value = 1");
               end
               96: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr1_inst.tdr[0:0], load value = 1");
               end
               97: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_tdr1_inst.tdr[0] ");
                  end
               end
               98: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_tdr2_inst.tdr[0] ");
                  end
               end
               99: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_tdr3_inst.tdr[0] ");
                  end
               end
               100: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_tdr4_inst.tdr[0] ");
                  end
               end
               101: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.sib, expected value = 1");
               end
               102: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.sib, expected value = 0");
               end
               103: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.sib, expected value = 0");
               end
               104: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.sib, expected value = 1");
               end
               105: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.sib, expected value = 1");
               end
               106: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr4_inst.tdr[0:0], expected value = 0");
               end
               107: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr3_inst.tdr[0:0], expected value = 0");
               end
               108: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr2_inst.tdr[0:0], expected value = 1");
               end
               109: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_tdr1_inst.tdr[0:0], expected value = 1");
               end
               110: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_sri_ctrl_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               111: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[13:0], load value = 10011110000111");
               end
               112: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[0] ");
                  end
               end
               113: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[1] ");
                  end
               end
               114: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[2] ");
                  end
               end
               115: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[3] ");
                  end
               end
               116: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[4] ");
                  end
               end
               117: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[5] ");
                  end
               end
               118: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[6] ");
                  end
               end
               119: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[7] ");
                  end
               end
               120: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[8] ");
                  end
               end
               121: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[9] ");
                  end
               end
               122: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[10] ");
                  end
               end
               123: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[11] ");
                  end
               end
               124: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[12] ");
                  end
               end
               125: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[13] ");
                  end
               end
               126: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_sri_ctrl_inst.tdr[13:0], expected value = 10011110000111");
               end
               127: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_edt_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               128: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_edt_intest_edt_tdr_inst.tdr[1:0], load value = 11");
               end
               129: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_edt_extest_edt_tdr_inst.tdr[1:0], load value = 00");
               end
               130: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_edt_intest_edt_tdr_inst.tdr[1:0], expected value = 11");
               end
               131: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_edt_extest_edt_tdr_inst.tdr[1:0], expected value = 00");
               end
               132: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_edt_extest_edt_tdr_inst.tdr[0] ");
                  end
               end
               133: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_edt_extest_edt_tdr_inst.tdr[1] ");
                  end
               end
               134: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_edt_intest_edt_tdr_inst.tdr[0] ");
                  end
               end
               135: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_edt_intest_edt_tdr_inst.tdr[1] ");
                  end
               end
               136: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_occ_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               137: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr_sib.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = scan_in");
               end
               138: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr_sib.sib, load value = 0");
               end
               139: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr_sib.sib ");
                  end
               end
               140: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr_sib.sib, expected value = 0");
               end
               141: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr_sib.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = from_scan_out");
               end
               142: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr[6:0], load value = 1111000");
               end
               143: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[0] ");
                  end
               end
               144: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[1] ");
                  end
               end
               145: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[2] ");
                  end
               end
               146: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[3] ");
                  end
               end
               147: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[4] ");
                  end
               end
               148: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[5] ");
                  end
               end
               149: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_occ_clk_inst.tdr[6] ");
                  end
               end
               150: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_occ_clk_inst.tdr[6:0], expected value = 1111000");
               end
               151: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_ssn_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               152: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.ijtag_so_mux, selection 3: config_sib_shift_reg, enable_shift_reg = 2'b11 -> ijtag_so_mux = enable_shift_reg");
               end
               153: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.streaming_through_ijtag_en_si_mux, selection 0: streaming_through_ijtag_en_si_mux_select = 1'b0 -> streaming_through_ijtag_en_si_mux = config_sib_shift_reg");
               end
               154: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_si_mux, selection 0: config_sib_shift_reg, enable_shift_reg = 2'b11 -> config_sib_si_mux = bus_out_shift_reg[0]");
               end
               155: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.enable_shift_reg ");
                  end
               end
               156: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[19:0], load value = 00111111111111111100");
               end
               157: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[19:0], load value = 11000011111111000000");
               end
               158: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_shift_reg, load value = 1");
               end
               159: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.enable_shift_reg, load value = 1");
               end
               160: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[19:0], expected value = 00111111111111111100");
               end
               161: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[19:0], expected value = 11000011111111000000");
               end
               162: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_shift_reg, expected value = 1");
               end
               163: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.enable_shift_reg, expected value = 1");
               end
               164: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_shift_reg ");
                  end
               end
               165: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[0] ");
                  end
               end
               166: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[1] ");
                  end
               end
               167: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[2] ");
                  end
               end
               168: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[3] ");
                  end
               end
               169: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[4] ");
                  end
               end
               170: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[5] ");
                  end
               end
               171: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[6] ");
                  end
               end
               172: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[7] ");
                  end
               end
               173: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[8] ");
                  end
               end
               174: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[9] ");
                  end
               end
               175: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[10] ");
                  end
               end
               176: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[11] ");
                  end
               end
               177: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[12] ");
                  end
               end
               178: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[13] ");
                  end
               end
               179: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[14] ");
                  end
               end
               180: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[15] ");
                  end
               end
               181: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[16] ");
                  end
               end
               182: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[17] ");
                  end
               end
               183: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[18] ");
                  end
               end
               184: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_out_shift_reg[19] ");
                  end
               end
               185: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[0] ");
                  end
               end
               186: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[1] ");
                  end
               end
               187: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[2] ");
                  end
               end
               188: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[3] ");
                  end
               end
               189: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[4] ");
                  end
               end
               190: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[5] ");
                  end
               end
               191: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[6] ");
                  end
               end
               192: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[7] ");
                  end
               end
               193: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[8] ");
                  end
               end
               194: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[9] ");
                  end
               end
               195: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[10] ");
                  end
               end
               196: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[11] ");
                  end
               end
               197: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[12] ");
                  end
               end
               198: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[13] ");
                  end
               end
               199: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[14] ");
                  end
               end
               200: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[15] ");
                  end
               end
               201: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[16] ");
                  end
               end
               202: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[17] ");
                  end
               end
               203: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[18] ");
                  end
               end
               204: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_in_shift_reg[19] ");
                  end
               end
               205: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.ijtag_so_mux, selection 1: config_sib_shift_reg, enable_shift_reg = 2'b00 -> ijtag_so_mux = enable_shift_reg");
               end
               206: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_si_mux, selection 1: config_sib_shift_reg, enable_shift_reg = 2'bxx -> config_sib_si_mux = ijtag_si");
               end
               207: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.ijtag_so_mux, selection 0: config_sib_shift_reg, enable_shift_reg = 2'b10 -> ijtag_so_mux = packet_width_is_less_than_two_bus_clock_shift_reg");
               end
               208: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_shift_reg, load value = 0");
               end
               209: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.enable_shift_reg, load value = 0");
               end
               210: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.streaming_through_ijtag_en_shift_reg, load value = 0");
               end
               211: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[30:0], load value = 1111111111111111111111111111100");
               end
               212: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.relative_initial_offset_enable_shift_reg, load value = 1");
               end
               213: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[4:0], load value = 11111");
               end
               214: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[8:0], load value = 111111111");
               end
               215: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.to_scan_in_bits_shift_reg[2:0], load value = 111");
               end
               216: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_bits_shift_reg[1:0], load value = 11");
               end
               217: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_le_strobe_en_shift_reg, load value = 1");
               end
               218: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[27:0], load value = 0000000000000011111111111111");
               end
               219: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[27:0], load value = 1111111111000000000000000000");
               end
               220: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[15:0], load value = 1111111111111111");
               end
               221: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.force_suppress_capture_shift_reg, load value = 1");
               end
               222: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[4:0], load value = 11111");
               end
               223: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_enable_shift_reg, load value = 0");
               end
               224: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_on_chip_compare_contribution_shift_reg, load value = 0");
               end
               225: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[7:0], load value = 00000000");
               end
               226: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[7:0], load value = 11000000");
               end
               227: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.loop_back_en_shift_reg, load value = 1");
               end
               228: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.capture_packets_shift_reg[2:0], load value = 111");
               end
               229: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.init_scan_load_used_shift_reg, load value = 1");
               end
               230: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_first_scan_load_masking_shift_reg, load value = 1");
               end
               231: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packets_per_capture_clock_minus_one_shift_reg[2:0], load value = 111");
               end
               232: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[3:0], load value = 1111");
               end
               233: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[3:0], load value = 0001");
               end
               234: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[3:0], load value = 0000");
               end
               235: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[3:0], load value = 1110");
               end
               236: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[5:0], load value = 011111");
               end
               237: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[5:0], load value = 111000");
               end
               238: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_width_is_less_than_two_bus_clock_shift_reg, load value = 1");
               end
               239: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.config_sib_shift_reg, expected value = 0");
               end
               240: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.enable_shift_reg, expected value = 0");
               end
               241: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.streaming_through_ijtag_en_shift_reg, expected value = 0");
               end
               242: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[30:0], expected value = 1111111111111111111111111111100");
               end
               243: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.relative_initial_offset_enable_shift_reg, expected value = 1");
               end
               244: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[4:0], expected value = 11111");
               end
               245: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[8:0], expected value = 111111111");
               end
               246: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.to_scan_in_bits_shift_reg[2:0], expected value = 111");
               end
               247: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_bits_shift_reg[1:0], expected value = 11");
               end
               248: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_le_strobe_en_shift_reg, expected value = 1");
               end
               249: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[27:0], expected value = 0000000000000011111111111111");
               end
               250: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[27:0], expected value = 1111111111000000000000000000");
               end
               251: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[15:0], expected value = 1111111111111111");
               end
               252: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.force_suppress_capture_shift_reg, expected value = 1");
               end
               253: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[4:0], expected value = 11111");
               end
               254: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_enable_shift_reg, expected value = 0");
               end
               255: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_on_chip_compare_contribution_shift_reg, expected value = 0");
               end
               256: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[7:0], expected value = 00000000");
               end
               257: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[7:0], expected value = 11000000");
               end
               258: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.loop_back_en_shift_reg, expected value = 1");
               end
               259: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.capture_packets_shift_reg[2:0], expected value = 111");
               end
               260: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.init_scan_load_used_shift_reg, expected value = 1");
               end
               261: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_first_scan_load_masking_shift_reg, expected value = 1");
               end
               262: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packets_per_capture_clock_minus_one_shift_reg[2:0], expected value = 111");
               end
               263: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[3:0], expected value = 1111");
               end
               264: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[3:0], expected value = 0001");
               end
               265: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[3:0], expected value = 0000");
               end
               266: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[3:0], expected value = 1110");
               end
               267: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[5:0], expected value = 011111");
               end
               268: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[5:0], expected value = 111000");
               end
               269: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_width_is_less_than_two_bus_clock_shift_reg, expected value = 1");
               end
               270: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_width_is_less_than_two_bus_clock_shift_reg ");
                  end
               end
               271: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[0] ");
                  end
               end
               272: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[1] ");
                  end
               end
               273: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[2] ");
                  end
               end
               274: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[3] ");
                  end
               end
               275: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[4] ");
                  end
               end
               276: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_capture_clock_low_width_shift_reg[5] ");
                  end
               end
               277: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[0] ");
                  end
               end
               278: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[1] ");
                  end
               end
               279: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[2] ");
                  end
               end
               280: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[3] ");
                  end
               end
               281: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[4] ");
                  end
               end
               282: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.min_shift_clock_low_width_shift_reg[5] ");
                  end
               end
               283: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[0] ");
                  end
               end
               284: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[1] ");
                  end
               end
               285: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[2] ");
                  end
               end
               286: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_launch_word_shift_reg[3] ");
                  end
               end
               287: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[0] ");
                  end
               end
               288: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[1] ");
                  end
               end
               289: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[2] ");
                  end
               end
               290: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.edt_update_falling_transition_words_shift_reg[3] ");
                  end
               end
               291: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[0] ");
                  end
               end
               292: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[1] ");
                  end
               end
               293: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[2] ");
                  end
               end
               294: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_launch_packet_shift_reg[3] ");
                  end
               end
               295: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[0] ");
                  end
               end
               296: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[1] ");
                  end
               end
               297: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[2] ");
                  end
               end
               298: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.scan_en_transition_packets_shift_reg[3] ");
                  end
               end
               299: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packets_per_capture_clock_minus_one_shift_reg[0] ");
                  end
               end
               300: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packets_per_capture_clock_minus_one_shift_reg[1] ");
                  end
               end
               301: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packets_per_capture_clock_minus_one_shift_reg[2] ");
                  end
               end
               302: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_first_scan_load_masking_shift_reg ");
                  end
               end
               303: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.init_scan_load_used_shift_reg ");
                  end
               end
               304: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.capture_packets_shift_reg[0] ");
                  end
               end
               305: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.capture_packets_shift_reg[1] ");
                  end
               end
               306: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.capture_packets_shift_reg[2] ");
                  end
               end
               307: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.loop_back_en_shift_reg ");
                  end
               end
               308: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[0] ");
                  end
               end
               309: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[1] ");
                  end
               end
               310: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[2] ");
                  end
               end
               311: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[3] ");
                  end
               end
               312: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[4] ");
                  end
               end
               313: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[5] ");
                  end
               end
               314: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[6] ");
                  end
               end
               315: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_shift_reg[7] ");
                  end
               end
               316: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[0] ");
                  end
               end
               317: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[1] ");
                  end
               end
               318: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[2] ");
                  end
               end
               319: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[3] ");
                  end
               end
               320: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[4] ");
                  end
               end
               321: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[5] ");
                  end
               end
               322: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[6] ");
                  end
               end
               323: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_group_count_shift_reg[7] ");
                  end
               end
               324: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.disable_on_chip_compare_contribution_shift_reg ");
                  end
               end
               325: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.on_chip_compare_enable_shift_reg ");
                  end
               end
               326: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[0] ");
                  end
               end
               327: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[1] ");
                  end
               end
               328: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[2] ");
                  end
               end
               329: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[3] ");
                  end
               end
               330: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_bit0_position_shift_reg[4] ");
                  end
               end
               331: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.force_suppress_capture_shift_reg ");
                  end
               end
               332: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[0] ");
                  end
               end
               333: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[1] ");
                  end
               end
               334: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[2] ");
                  end
               end
               335: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[3] ");
                  end
               end
               336: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[4] ");
                  end
               end
               337: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[5] ");
                  end
               end
               338: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[6] ");
                  end
               end
               339: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[7] ");
                  end
               end
               340: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[8] ");
                  end
               end
               341: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[9] ");
                  end
               end
               342: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[10] ");
                  end
               end
               343: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[11] ");
                  end
               end
               344: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[12] ");
                  end
               end
               345: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[13] ");
                  end
               end
               346: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[14] ");
                  end
               end
               347: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.packet_size_shift_reg[15] ");
                  end
               end
               348: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[0] ");
                  end
               end
               349: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[1] ");
                  end
               end
               350: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[2] ");
                  end
               end
               351: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[3] ");
                  end
               end
               352: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[4] ");
                  end
               end
               353: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[5] ");
                  end
               end
               354: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[6] ");
                  end
               end
               355: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[7] ");
                  end
               end
               356: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[8] ");
                  end
               end
               357: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[9] ");
                  end
               end
               358: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[10] ");
                  end
               end
               359: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[11] ");
                  end
               end
               360: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[12] ");
                  end
               end
               361: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[13] ");
                  end
               end
               362: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[14] ");
                  end
               end
               363: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[15] ");
                  end
               end
               364: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[16] ");
                  end
               end
               365: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[17] ");
                  end
               end
               366: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[18] ");
                  end
               end
               367: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[19] ");
                  end
               end
               368: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[20] ");
                  end
               end
               369: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[21] ");
                  end
               end
               370: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[22] ");
                  end
               end
               371: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[23] ");
                  end
               end
               372: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[24] ");
                  end
               end
               373: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[25] ");
                  end
               end
               374: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[26] ");
                  end
               end
               375: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.extra_shift_packets_shift_reg[27] ");
                  end
               end
               376: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[0] ");
                  end
               end
               377: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[1] ");
                  end
               end
               378: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[2] ");
                  end
               end
               379: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[3] ");
                  end
               end
               380: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[4] ");
                  end
               end
               381: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[5] ");
                  end
               end
               382: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[6] ");
                  end
               end
               383: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[7] ");
                  end
               end
               384: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[8] ");
                  end
               end
               385: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[9] ");
                  end
               end
               386: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[10] ");
                  end
               end
               387: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[11] ");
                  end
               end
               388: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[12] ");
                  end
               end
               389: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[13] ");
                  end
               end
               390: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[14] ");
                  end
               end
               391: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[15] ");
                  end
               end
               392: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[16] ");
                  end
               end
               393: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[17] ");
                  end
               end
               394: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[18] ");
                  end
               end
               395: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[19] ");
                  end
               end
               396: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[20] ");
                  end
               end
               397: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[21] ");
                  end
               end
               398: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[22] ");
                  end
               end
               399: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[23] ");
                  end
               end
               400: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[24] ");
                  end
               end
               401: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[25] ");
                  end
               end
               402: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[26] ");
                  end
               end
               403: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.total_shift_cnt_minus_one_shift_reg[27] ");
                  end
               end
               404: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_le_strobe_en_shift_reg ");
                  end
               end
               405: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_bits_shift_reg[0] ");
                  end
               end
               406: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.from_scan_out_bits_shift_reg[1] ");
                  end
               end
               407: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.to_scan_in_bits_shift_reg[0] ");
                  end
               end
               408: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.to_scan_in_bits_shift_reg[1] ");
                  end
               end
               409: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.to_scan_in_bits_shift_reg[2] ");
                  end
               end
               410: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[0] ");
                  end
               end
               411: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[1] ");
                  end
               end
               412: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[2] ");
                  end
               end
               413: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[3] ");
                  end
               end
               414: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[4] ");
                  end
               end
               415: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[5] ");
                  end
               end
               416: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[6] ");
                  end
               end
               417: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[7] ");
                  end
               end
               418: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bits_per_packet_shift_reg[8] ");
                  end
               end
               419: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[0] ");
                  end
               end
               420: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[1] ");
                  end
               end
               421: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[2] ");
                  end
               end
               422: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[3] ");
                  end
               end
               423: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.bus_width_shift_reg[4] ");
                  end
               end
               424: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.relative_initial_offset_enable_shift_reg ");
                  end
               end
               425: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[0] ");
                  end
               end
               426: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[1] ");
                  end
               end
               427: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[2] ");
                  end
               end
               428: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[3] ");
                  end
               end
               429: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[4] ");
                  end
               end
               430: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[5] ");
                  end
               end
               431: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[6] ");
                  end
               end
               432: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[7] ");
                  end
               end
               433: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[8] ");
                  end
               end
               434: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[9] ");
                  end
               end
               435: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[10] ");
                  end
               end
               436: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[11] ");
                  end
               end
               437: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[12] ");
                  end
               end
               438: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[13] ");
                  end
               end
               439: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[14] ");
                  end
               end
               440: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[15] ");
                  end
               end
               441: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[16] ");
                  end
               end
               442: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[17] ");
                  end
               end
               443: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[18] ");
                  end
               end
               444: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[19] ");
                  end
               end
               445: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[20] ");
                  end
               end
               446: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[21] ");
                  end
               end
               447: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[22] ");
                  end
               end
               448: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[23] ");
                  end
               end
               449: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[24] ");
                  end
               end
               450: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[25] ");
                  end
               end
               451: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[26] ");
                  end
               end
               452: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[27] ");
                  end
               end
               453: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[28] ");
                  end
               end
               454: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[29] ");
                  end
               end
               455: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.initial_offset_shift_reg[30] ");
                  end
               end
               456: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_ssn_scan_host_ssh_inst.inner.streaming_through_ijtag_en_shift_reg ");
                  end
               end
               457: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_intest_edt_scan_bi_sol_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               458: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_intest_edt_scan_bi_sol_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               459: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_intest_edt_scan_bi_sol_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               460: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[20:0], load value = 110000000011111111111");
               end
               461: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[17:0], load value = 110011110000111111");
               end
               462: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[20:0], expected value = 110000000011111111111");
               end
               463: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[17:0], expected value = 110011110000111111");
               end
               464: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[0] ");
                  end
               end
               465: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[1] ");
                  end
               end
               466: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[2] ");
                  end
               end
               467: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[3] ");
                  end
               end
               468: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[4] ");
                  end
               end
               469: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[5] ");
                  end
               end
               470: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[6] ");
                  end
               end
               471: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[7] ");
                  end
               end
               472: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[8] ");
                  end
               end
               473: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[9] ");
                  end
               end
               474: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[10] ");
                  end
               end
               475: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[11] ");
                  end
               end
               476: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[12] ");
                  end
               end
               477: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[13] ");
                  end
               end
               478: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[14] ");
                  end
               end
               479: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[15] ");
                  end
               end
               480: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[16] ");
                  end
               end
               481: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_status_inst.tdr[17] ");
                  end
               end
               482: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[0] ");
                  end
               end
               483: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[1] ");
                  end
               end
               484: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[2] ");
                  end
               end
               485: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[3] ");
                  end
               end
               486: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[4] ");
                  end
               end
               487: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[5] ");
                  end
               end
               488: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[6] ");
                  end
               end
               489: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[7] ");
                  end
               end
               490: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[8] ");
                  end
               end
               491: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[9] ");
                  end
               end
               492: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[10] ");
                  end
               end
               493: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[11] ");
                  end
               end
               494: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[12] ");
                  end
               end
               495: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[13] ");
                  end
               end
               496: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[14] ");
                  end
               end
               497: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[15] ");
                  end
               end
               498: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[16] ");
                  end
               end
               499: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[17] ");
                  end
               end
               500: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[18] ");
                  end
               end
               501: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[19] ");
                  end
               end
               502: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_intest_edt_scan_bi_sol_control_inst.tdr[20] ");
                  end
               end
               503: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_sib_extest_edt_scan_bi_sol_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               504: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_extest_edt_scan_bi_sol_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               505: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_scanmux_extest_edt_scan_bi_sol_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               506: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[19:0], load value = 11000000001111111111");
               end
               507: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[16:0], load value = 10011110000111111");
               end
               508: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[19:0], expected value = 11000000001111111111");
               end
               509: begin
                  $display($realtime, "ns:   firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[16:0], expected value = 10011110000111111");
               end
               510: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[0] ");
                  end
               end
               511: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[1] ");
                  end
               end
               512: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[2] ");
                  end
               end
               513: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[3] ");
                  end
               end
               514: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[4] ");
                  end
               end
               515: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[5] ");
                  end
               end
               516: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[6] ");
                  end
               end
               517: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[7] ");
                  end
               end
               518: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[8] ");
                  end
               end
               519: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[9] ");
                  end
               end
               520: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[10] ");
                  end
               end
               521: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[11] ");
                  end
               end
               522: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[12] ");
                  end
               end
               523: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[13] ");
                  end
               end
               524: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[14] ");
                  end
               end
               525: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[15] ");
                  end
               end
               526: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_status_inst.tdr[16] ");
                  end
               end
               527: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[0] ");
                  end
               end
               528: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[1] ");
                  end
               end
               529: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[2] ");
                  end
               end
               530: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[3] ");
                  end
               end
               531: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[4] ");
                  end
               end
               532: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[5] ");
                  end
               end
               533: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[6] ");
                  end
               end
               534: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[7] ");
                  end
               end
               535: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[8] ");
                  end
               end
               536: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[9] ");
                  end
               end
               537: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[10] ");
                  end
               end
               538: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[11] ");
                  end
               end
               539: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[12] ");
                  end
               end
               540: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[13] ");
                  end
               end
               541: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[14] ");
                  end
               end
               542: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[15] ");
                  end
               end
               543: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[16] ");
                  end
               end
               544: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[17] ");
                  end
               end
               545: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[18] ");
                  end
               end
               546: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate2_tessent_tdr_extest_edt_scan_bi_sol_control_inst.tdr[19] ");
                  end
               end
               547: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_sti_inst.scan_in_mux, selection 0: sib, ltest_en = 2'b10 -> scan_in_mux = ijtag_from_so");
               end
               548: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_sti_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               549: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_sti_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               550: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_mbist_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               551: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_mbist_inst.sib, load value = 0");
               end
               552: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_sti_ctrl_inst.tdr[0:0], load value = 0");
               end
               553: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_mbist_inst.sib ");
                  end
               end
               554: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_mbist_inst.sib, expected value = 0");
               end
               555: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_sti_ctrl_inst.tdr[0:0], expected value = 0");
               end
               556: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_sti_ctrl_inst.tdr[0] ");
                  end
               end
               557: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_mbist_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               558: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.DiagnosisReadyScanMux, selection 0: sib = 1'b0 -> DiagnosisReadyScanMux = ijtag_si");
               end
               559: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ctl_sib_mux_inst, selection 0: ctl_group_sib = 1'b0 -> ctl_sib_mux_inst = tdr_bypass_sib_inst");
               end
               560: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_mux_inst, selection 0: tdr_bypass_sib_inst = 1'b0 -> tdr_bypass_sib_mux_inst = si");
               end
               561: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_inst, load value = 1");
               end
               562: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ctl_group_sib, load value = 1");
               end
               563: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.sib, load value = 1");
               end
               564: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ctl_group_sib ");
                  end
               end
               565: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_inst ");
                  end
               end
               566: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_inst, expected value = 1");
               end
               567: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ctl_group_sib, expected value = 1");
               end
               568: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.sib, expected value = 1");
               end
               569: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.sib ");
                  end
               end
               570: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.DiagnosisReadyScanMux, selection 1: sib = 1'b1 -> DiagnosisReadyScanMux = tdr");
               end
               571: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.tdr, load value = 1");
               end
               572: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.tdr ");
                  end
               end
               573: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_diagnosis_ready_inst.tdr, expected value = 1");
               end
               574: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ctl_sib_mux_inst, selection 1: ctl_group_sib = 1'b1 -> ctl_sib_mux_inst = mbist_go_0");
               end
               575: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.fromBistMux_0, selection 1: bistEn_int[0], BIST_SETUP_tdr[1], ChainBypassMode = 3'bxxx -> fromBistMux_0 = tdr_bypass_sib_inst");
               end
               576: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_inst, load value = 0");
               end
               577: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_done_0, load value = 1");
               end
               578: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_go_0, load value = 1");
               end
               579: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_inst, expected value = 0");
               end
               580: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_done_0, expected value = 1");
               end
               581: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_go_0, expected value = 1");
               end
               582: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_go_0 ");
                  end
               end
               583: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.mbist_done_0 ");
                  end
               end
               584: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.tdr_bypass_sib_mux_inst, selection 1: tdr_bypass_sib_inst = 1'b1 -> tdr_bypass_sib_mux_inst = ENABLE_MEM_RESET_tdr");
               end
               585: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SETUP_tdr[2:0], load value = 000");
               end
               586: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.TCK_MODE_tdr, load value = 0");
               end
               587: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHAIN_BYPASS_EN_tdr, load value = 0");
               end
               588: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.INCLUDE_MEM_RESULTS_REG_tdr, load value = 0");
               end
               589: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE1_tdr, load value = 1");
               end
               590: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE0_tdr, load value = 1");
               end
               591: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ASYNC_RESET_tdr, load value = 1");
               end
               592: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHECK_REPAIR_NEEDED_tdr, load value = 1");
               end
               593: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.PRESERVE_FUSE_REGISTER_tdr, load value = 1");
               end
               594: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_DIAG_EN_tdr, load value = 1");
               end
               595: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIRA_EN_tdr, load value = 1");
               end
               596: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.MEM_ARRAY_DUMP_MODE_tdr, load value = 1");
               end
               597: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE1_tdr, load value = 0");
               end
               598: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE0_tdr, load value = 0");
               end
               599: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SELECT_TEST_DATA_tdr, load value = 0");
               end
               600: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.REDUCED_ADDRESS_COUNT_tdr, load value = 0");
               end
               601: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ENABLE_MEM_RESET_tdr, load value = 1");
               end
               602: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SETUP_tdr[2:0], expected value = 000");
               end
               603: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.TCK_MODE_tdr, expected value = 0");
               end
               604: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHAIN_BYPASS_EN_tdr, expected value = 0");
               end
               605: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.INCLUDE_MEM_RESULTS_REG_tdr, expected value = 0");
               end
               606: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE1_tdr, expected value = 1");
               end
               607: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE0_tdr, expected value = 1");
               end
               608: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ASYNC_RESET_tdr, expected value = 1");
               end
               609: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHECK_REPAIR_NEEDED_tdr, expected value = 1");
               end
               610: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.PRESERVE_FUSE_REGISTER_tdr, expected value = 1");
               end
               611: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_DIAG_EN_tdr, expected value = 1");
               end
               612: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIRA_EN_tdr, expected value = 1");
               end
               613: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.MEM_ARRAY_DUMP_MODE_tdr, expected value = 1");
               end
               614: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE1_tdr, expected value = 0");
               end
               615: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE0_tdr, expected value = 0");
               end
               616: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SELECT_TEST_DATA_tdr, expected value = 0");
               end
               617: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.REDUCED_ADDRESS_COUNT_tdr, expected value = 0");
               end
               618: begin
                  $display($realtime, "ns:   ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ENABLE_MEM_RESET_tdr, expected value = 1");
               end
               619: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.ENABLE_MEM_RESET_tdr ");
                  end
               end
               620: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.REDUCED_ADDRESS_COUNT_tdr ");
                  end
               end
               621: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SELECT_TEST_DATA_tdr ");
                  end
               end
               622: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE0_tdr ");
                  end
               end
               623: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ALGO_MODE1_tdr ");
                  end
               end
               624: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.MEM_ARRAY_DUMP_MODE_tdr ");
                  end
               end
               625: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIRA_EN_tdr ");
                  end
               end
               626: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_DIAG_EN_tdr ");
                  end
               end
               627: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.PRESERVE_FUSE_REGISTER_tdr ");
                  end
               end
               628: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHECK_REPAIR_NEEDED_tdr ");
                  end
               end
               629: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_ASYNC_RESET_tdr ");
                  end
               end
               630: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE0_tdr ");
                  end
               end
               631: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.FL_CNT_MODE1_tdr ");
                  end
               end
               632: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.INCLUDE_MEM_RESULTS_REG_tdr ");
                  end
               end
               633: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.CHAIN_BYPASS_EN_tdr ");
                  end
               end
               634: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.TCK_MODE_tdr ");
                  end
               end
               635: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SETUP_tdr[0] ");
                  end
               end
               636: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SETUP_tdr[1] ");
                  end
               end
               637: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_firebird7_in_gate1_tessent_mbist_bap_inst.BIST_SETUP_tdr[2] ");
                  end
               end
               638: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               639: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_red_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               640: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_orange_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               641: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_insysbist_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               642: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_green_inst.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = ijtag_si");
               end
               643: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_green_inst.sib, load value = 1");
               end
               644: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_insysbist_inst.sib, load value = 1");
               end
               645: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_orange_inst.sib, load value = 1");
               end
               646: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_red_inst.sib, load value = 0");
               end
               647: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_spare_red_inst.sib ");
                  end
               end
               648: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_spare_orange_inst.sib ");
                  end
               end
               649: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_spare_insysbist_inst.sib ");
                  end
               end
               650: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_sib_spare_green_inst.sib ");
                  end
               end
               651: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_green_inst.sib, expected value = 1");
               end
               652: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_insysbist_inst.sib, expected value = 1");
               end
               653: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_orange_inst.sib, expected value = 1");
               end
               654: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_red_inst.sib, expected value = 0");
               end
               655: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_red_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               656: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_red_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               657: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_red_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               658: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[7:0], load value = 11110000");
               end
               659: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[7:0], expected value = 11110000");
               end
               660: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[0] ");
                  end
               end
               661: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[1] ");
                  end
               end
               662: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[2] ");
                  end
               end
               663: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[3] ");
                  end
               end
               664: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[4] ");
                  end
               end
               665: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[5] ");
                  end
               end
               666: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[6] ");
                  end
               end
               667: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_red_tdr_inst.tdr[7] ");
                  end
               end
               668: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_orange_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               669: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_orange_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               670: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_orange_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               671: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[7:0], load value = 11100001");
               end
               672: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[7:0], expected value = 11100001");
               end
               673: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[0] ");
                  end
               end
               674: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[1] ");
                  end
               end
               675: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[2] ");
                  end
               end
               676: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[3] ");
                  end
               end
               677: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[4] ");
                  end
               end
               678: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[5] ");
                  end
               end
               679: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[6] ");
                  end
               end
               680: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_orange_tdr_inst.tdr[7] ");
                  end
               end
               681: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_insysbist_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               682: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_insysbist_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               683: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_spare_insysbist_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               684: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[7:0], load value = 11000011");
               end
               685: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[7:0], expected value = 11000011");
               end
               686: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[0] ");
                  end
               end
               687: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[1] ");
                  end
               end
               688: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[2] ");
                  end
               end
               689: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[3] ");
                  end
               end
               690: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[4] ");
                  end
               end
               691: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[5] ");
                  end
               end
               692: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[6] ");
                  end
               end
               693: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_insysbist_tdr_inst.tdr[7] ");
                  end
               end
               694: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_spare_green_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               695: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[7:0], load value = 10000111");
               end
               696: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[7:0], expected value = 10000111");
               end
               697: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[0] ");
                  end
               end
               698: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[1] ");
                  end
               end
               699: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[2] ");
                  end
               end
               700: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[3] ");
                  end
               end
               701: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[4] ");
                  end
               end
               702: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[5] ");
                  end
               end
               703: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[6] ");
                  end
               end
               704: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = firebird7_in_gate1_tessent_tdr_spare_green_tdr_inst.tdr[7] ");
                  end
               end
               705: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_upm_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               706: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_upm_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               707: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_upm_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               708: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               709: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               710: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               711: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_CBB.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               712: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               713: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               714: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               715: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               716: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               717: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               718: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               719: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_CBB.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               720: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               721: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               722: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               723: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.scan_in_mux, selection 0: sib = 1'b0 -> scan_in_mux = si");
               end
               724: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.sib[0:0], load value = 1");
               end
               725: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 1");
               end
               726: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 1");
               end
               727: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 1");
               end
               728: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_CBB.sib[0:0], load value = 1");
               end
               729: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 1");
               end
               730: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 1");
               end
               731: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 1");
               end
               732: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.sib[0:0], load value = 0");
               end
               733: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 0");
               end
               734: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 0");
               end
               735: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 0");
               end
               736: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_CBB.sib[0:0], load value = 1");
               end
               737: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 1");
               end
               738: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 1");
               end
               739: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 1");
               end
               740: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.sib[0:0], expected value = 1");
               end
               741: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 1");
               end
               742: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 1");
               end
               743: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 1");
               end
               744: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_CBB.sib[0:0], expected value = 1");
               end
               745: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 1");
               end
               746: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 1");
               end
               747: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 1");
               end
               748: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.sib[0:0], expected value = 0");
               end
               749: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 0");
               end
               750: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 0");
               end
               751: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 0");
               end
               752: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_CBB.sib[0:0], expected value = 1");
               end
               753: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 1");
               end
               754: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 1");
               end
               755: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 1");
               end
               756: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.SIB_UPM_STATUS.sib[0] ");
                  end
               end
               757: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.SIB_COUNTER_RESULT.sib[0] ");
                  end
               end
               758: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.SIB_COUNTER_CTRL.sib[0] ");
                  end
               end
               759: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.SIB_CBB.sib[0] ");
                  end
               end
               760: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.SIB_UPM_STATUS.sib[0] ");
                  end
               end
               761: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.SIB_COUNTER_RESULT.sib[0] ");
                  end
               end
               762: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.SIB_COUNTER_CTRL.sib[0] ");
                  end
               end
               763: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.SIB_CBB.sib[0] ");
                  end
               end
               764: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.SIB_UPM_STATUS.sib[0] ");
                  end
               end
               765: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.SIB_COUNTER_RESULT.sib[0] ");
                  end
               end
               766: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.SIB_COUNTER_CTRL.sib[0] ");
                  end
               end
               767: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.SIB_CBB.sib[0] ");
                  end
               end
               768: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.SIB_UPM_STATUS.sib[0] ");
                  end
               end
               769: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.SIB_COUNTER_RESULT.sib[0] ");
                  end
               end
               770: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.SIB_COUNTER_CTRL.sib[0] ");
                  end
               end
               771: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.SIB_CBB.sib[0] ");
                  end
               end
               772: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               773: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.sib[0:0], load value = 0");
               end
               774: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.sib[0:0], load value = 1");
               end
               775: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 1");
               end
               776: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 1");
               end
               777: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 1");
               end
               778: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.UPM_STATUS_reg.DR[24:0], load value = 1110000111111110000000011");
               end
               779: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.sib[0:0], expected value = 0");
               end
               780: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.sib[0:0], expected value = 1");
               end
               781: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 1");
               end
               782: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 1");
               end
               783: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 1");
               end
               784: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.UPM_STATUS_reg.DR[24:0], expected value = 1110000111111110000000011");
               end
               785: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[0] ");
                  end
               end
               786: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[1] ");
                  end
               end
               787: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[2] ");
                  end
               end
               788: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[3] ");
                  end
               end
               789: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[4] ");
                  end
               end
               790: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[5] ");
                  end
               end
               791: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[6] ");
                  end
               end
               792: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[7] ");
                  end
               end
               793: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[8] ");
                  end
               end
               794: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[9] ");
                  end
               end
               795: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[10] ");
                  end
               end
               796: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[11] ");
                  end
               end
               797: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[12] ");
                  end
               end
               798: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[13] ");
                  end
               end
               799: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[14] ");
                  end
               end
               800: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[15] ");
                  end
               end
               801: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[16] ");
                  end
               end
               802: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[17] ");
                  end
               end
               803: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[18] ");
                  end
               end
               804: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[19] ");
                  end
               end
               805: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[20] ");
                  end
               end
               806: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[21] ");
                  end
               end
               807: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[22] ");
                  end
               end
               808: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[23] ");
                  end
               end
               809: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.UPM_STATUS_reg.DR[24] ");
                  end
               end
               810: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               811: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 0");
               end
               812: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[20:0], load value = 110000111111110000000");
               end
               813: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 0");
               end
               814: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[20:0], expected value = 110000111111110000000");
               end
               815: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[0] ");
                  end
               end
               816: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[1] ");
                  end
               end
               817: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[2] ");
                  end
               end
               818: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[3] ");
                  end
               end
               819: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[4] ");
                  end
               end
               820: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[5] ");
                  end
               end
               821: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[6] ");
                  end
               end
               822: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[7] ");
                  end
               end
               823: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[8] ");
                  end
               end
               824: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[9] ");
                  end
               end
               825: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[10] ");
                  end
               end
               826: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[11] ");
                  end
               end
               827: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[12] ");
                  end
               end
               828: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[13] ");
                  end
               end
               829: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[14] ");
                  end
               end
               830: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[15] ");
                  end
               end
               831: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[16] ");
                  end
               end
               832: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[17] ");
                  end
               end
               833: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[18] ");
                  end
               end
               834: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[19] ");
                  end
               end
               835: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_RESULT_reg.DR[20] ");
                  end
               end
               836: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               837: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.sib[0:0], load value = 0");
               end
               838: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[25:0], load value = 10000111111110000000011111");
               end
               839: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.sib[0:0], expected value = 0");
               end
               840: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[25:0], expected value = 10000111111110000000011111");
               end
               841: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[0] ");
                  end
               end
               842: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[1] ");
                  end
               end
               843: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[2] ");
                  end
               end
               844: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[3] ");
                  end
               end
               845: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[4] ");
                  end
               end
               846: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[5] ");
                  end
               end
               847: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[6] ");
                  end
               end
               848: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[7] ");
                  end
               end
               849: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[8] ");
                  end
               end
               850: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[9] ");
                  end
               end
               851: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[10] ");
                  end
               end
               852: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[11] ");
                  end
               end
               853: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[12] ");
                  end
               end
               854: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[13] ");
                  end
               end
               855: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[14] ");
                  end
               end
               856: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[15] ");
                  end
               end
               857: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[16] ");
                  end
               end
               858: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[17] ");
                  end
               end
               859: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[18] ");
                  end
               end
               860: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[19] ");
                  end
               end
               861: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[20] ");
                  end
               end
               862: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[21] ");
                  end
               end
               863: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[22] ");
                  end
               end
               864: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[23] ");
                  end
               end
               865: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[24] ");
                  end
               end
               866: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.COUNTER_CTRL_reg.DR[25] ");
                  end
               end
               867: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.SIB_CBB.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               868: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.sib[0:0], load value = 0");
               end
               869: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.sib[0:0], load value = 0");
               end
               870: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.CBB_reg.DR[27:0], load value = 0000111111110000000011111111");
               end
               871: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.sib[0:0], expected value = 0");
               end
               872: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.sib[0:0], expected value = 0");
               end
               873: begin
                  $display($realtime, "ns:   u_upm_0.upm_inst.CBB_reg.DR[27:0], expected value = 0000111111110000000011111111");
               end
               874: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[0] ");
                  end
               end
               875: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[1] ");
                  end
               end
               876: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[2] ");
                  end
               end
               877: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[3] ");
                  end
               end
               878: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[4] ");
                  end
               end
               879: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[5] ");
                  end
               end
               880: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[6] ");
                  end
               end
               881: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[7] ");
                  end
               end
               882: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[8] ");
                  end
               end
               883: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[9] ");
                  end
               end
               884: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[10] ");
                  end
               end
               885: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[11] ");
                  end
               end
               886: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[12] ");
                  end
               end
               887: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[13] ");
                  end
               end
               888: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[14] ");
                  end
               end
               889: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[15] ");
                  end
               end
               890: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[16] ");
                  end
               end
               891: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[17] ");
                  end
               end
               892: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[18] ");
                  end
               end
               893: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[19] ");
                  end
               end
               894: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[20] ");
                  end
               end
               895: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[21] ");
                  end
               end
               896: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[22] ");
                  end
               end
               897: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[23] ");
                  end
               end
               898: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[24] ");
                  end
               end
               899: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[25] ");
                  end
               end
               900: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[26] ");
                  end
               end
               901: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_0.upm_inst.CBB_reg.DR[27] ");
                  end
               end
               902: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               903: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.UPM_STATUS_reg.DR[24:0], load value = 0001111111100000000111111");
               end
               904: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.UPM_STATUS_reg.DR[24:0], expected value = 0001111111100000000111111");
               end
               905: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[0] ");
                  end
               end
               906: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[1] ");
                  end
               end
               907: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[2] ");
                  end
               end
               908: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[3] ");
                  end
               end
               909: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[4] ");
                  end
               end
               910: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[5] ");
                  end
               end
               911: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[6] ");
                  end
               end
               912: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[7] ");
                  end
               end
               913: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[8] ");
                  end
               end
               914: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[9] ");
                  end
               end
               915: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[10] ");
                  end
               end
               916: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[11] ");
                  end
               end
               917: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[12] ");
                  end
               end
               918: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[13] ");
                  end
               end
               919: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[14] ");
                  end
               end
               920: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[15] ");
                  end
               end
               921: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[16] ");
                  end
               end
               922: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[17] ");
                  end
               end
               923: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[18] ");
                  end
               end
               924: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[19] ");
                  end
               end
               925: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[20] ");
                  end
               end
               926: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[21] ");
                  end
               end
               927: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[22] ");
                  end
               end
               928: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[23] ");
                  end
               end
               929: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.UPM_STATUS_reg.DR[24] ");
                  end
               end
               930: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               931: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[20:0], load value = 001111111100000000111");
               end
               932: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[20:0], expected value = 001111111100000000111");
               end
               933: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[0] ");
                  end
               end
               934: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[1] ");
                  end
               end
               935: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[2] ");
                  end
               end
               936: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[3] ");
                  end
               end
               937: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[4] ");
                  end
               end
               938: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[5] ");
                  end
               end
               939: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[6] ");
                  end
               end
               940: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[7] ");
                  end
               end
               941: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[8] ");
                  end
               end
               942: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[9] ");
                  end
               end
               943: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[10] ");
                  end
               end
               944: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[11] ");
                  end
               end
               945: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[12] ");
                  end
               end
               946: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[13] ");
                  end
               end
               947: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[14] ");
                  end
               end
               948: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[15] ");
                  end
               end
               949: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[16] ");
                  end
               end
               950: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[17] ");
                  end
               end
               951: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[18] ");
                  end
               end
               952: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[19] ");
                  end
               end
               953: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_RESULT_reg.DR[20] ");
                  end
               end
               954: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               955: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[25:0], load value = 01111111100000000111111111");
               end
               956: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[25:0], expected value = 01111111100000000111111111");
               end
               957: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[0] ");
                  end
               end
               958: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[1] ");
                  end
               end
               959: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[2] ");
                  end
               end
               960: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[3] ");
                  end
               end
               961: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[4] ");
                  end
               end
               962: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[5] ");
                  end
               end
               963: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[6] ");
                  end
               end
               964: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[7] ");
                  end
               end
               965: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[8] ");
                  end
               end
               966: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[9] ");
                  end
               end
               967: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[10] ");
                  end
               end
               968: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[11] ");
                  end
               end
               969: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[12] ");
                  end
               end
               970: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[13] ");
                  end
               end
               971: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[14] ");
                  end
               end
               972: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[15] ");
                  end
               end
               973: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[16] ");
                  end
               end
               974: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[17] ");
                  end
               end
               975: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[18] ");
                  end
               end
               976: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[19] ");
                  end
               end
               977: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[20] ");
                  end
               end
               978: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[21] ");
                  end
               end
               979: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[22] ");
                  end
               end
               980: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[23] ");
                  end
               end
               981: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[24] ");
                  end
               end
               982: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.COUNTER_CTRL_reg.DR[25] ");
                  end
               end
               983: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.SIB_CBB.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               984: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.CBB_reg.DR[27:0], load value = 1111111100000000111111111111");
               end
               985: begin
                  $display($realtime, "ns:   u_upm_1.upm_inst.CBB_reg.DR[27:0], expected value = 1111111100000000111111111111");
               end
               986: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[0] ");
                  end
               end
               987: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[1] ");
                  end
               end
               988: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[2] ");
                  end
               end
               989: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[3] ");
                  end
               end
               990: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[4] ");
                  end
               end
               991: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[5] ");
                  end
               end
               992: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[6] ");
                  end
               end
               993: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[7] ");
                  end
               end
               994: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[8] ");
                  end
               end
               995: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[9] ");
                  end
               end
               996: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[10] ");
                  end
               end
               997: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[11] ");
                  end
               end
               998: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[12] ");
                  end
               end
               999: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[13] ");
                  end
               end
               1000: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[14] ");
                  end
               end
               1001: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[15] ");
                  end
               end
               1002: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[16] ");
                  end
               end
               1003: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[17] ");
                  end
               end
               1004: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[18] ");
                  end
               end
               1005: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[19] ");
                  end
               end
               1006: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[20] ");
                  end
               end
               1007: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[21] ");
                  end
               end
               1008: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[22] ");
                  end
               end
               1009: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[23] ");
                  end
               end
               1010: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[24] ");
                  end
               end
               1011: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[25] ");
                  end
               end
               1012: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[26] ");
                  end
               end
               1013: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_1.upm_inst.CBB_reg.DR[27] ");
                  end
               end
               1014: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1015: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.UPM_STATUS_reg.DR[24:0], load value = 1111111000000001111111111");
               end
               1016: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.UPM_STATUS_reg.DR[24:0], expected value = 1111111000000001111111111");
               end
               1017: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[0] ");
                  end
               end
               1018: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[1] ");
                  end
               end
               1019: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[2] ");
                  end
               end
               1020: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[3] ");
                  end
               end
               1021: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[4] ");
                  end
               end
               1022: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[5] ");
                  end
               end
               1023: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[6] ");
                  end
               end
               1024: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[7] ");
                  end
               end
               1025: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[8] ");
                  end
               end
               1026: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[9] ");
                  end
               end
               1027: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[10] ");
                  end
               end
               1028: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[11] ");
                  end
               end
               1029: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[12] ");
                  end
               end
               1030: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[13] ");
                  end
               end
               1031: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[14] ");
                  end
               end
               1032: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[15] ");
                  end
               end
               1033: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[16] ");
                  end
               end
               1034: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[17] ");
                  end
               end
               1035: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[18] ");
                  end
               end
               1036: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[19] ");
                  end
               end
               1037: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[20] ");
                  end
               end
               1038: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[21] ");
                  end
               end
               1039: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[22] ");
                  end
               end
               1040: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[23] ");
                  end
               end
               1041: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.UPM_STATUS_reg.DR[24] ");
                  end
               end
               1042: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1043: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[20:0], load value = 111111000000001111111");
               end
               1044: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[20:0], expected value = 111111000000001111111");
               end
               1045: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[0] ");
                  end
               end
               1046: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[1] ");
                  end
               end
               1047: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[2] ");
                  end
               end
               1048: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[3] ");
                  end
               end
               1049: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[4] ");
                  end
               end
               1050: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[5] ");
                  end
               end
               1051: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[6] ");
                  end
               end
               1052: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[7] ");
                  end
               end
               1053: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[8] ");
                  end
               end
               1054: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[9] ");
                  end
               end
               1055: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[10] ");
                  end
               end
               1056: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[11] ");
                  end
               end
               1057: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[12] ");
                  end
               end
               1058: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[13] ");
                  end
               end
               1059: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[14] ");
                  end
               end
               1060: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[15] ");
                  end
               end
               1061: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[16] ");
                  end
               end
               1062: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[17] ");
                  end
               end
               1063: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[18] ");
                  end
               end
               1064: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[19] ");
                  end
               end
               1065: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_RESULT_reg.DR[20] ");
                  end
               end
               1066: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1067: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[25:0], load value = 11111000000001111111111111");
               end
               1068: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[25:0], expected value = 11111000000001111111111111");
               end
               1069: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[0] ");
                  end
               end
               1070: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[1] ");
                  end
               end
               1071: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[2] ");
                  end
               end
               1072: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[3] ");
                  end
               end
               1073: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[4] ");
                  end
               end
               1074: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[5] ");
                  end
               end
               1075: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[6] ");
                  end
               end
               1076: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[7] ");
                  end
               end
               1077: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[8] ");
                  end
               end
               1078: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[9] ");
                  end
               end
               1079: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[10] ");
                  end
               end
               1080: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[11] ");
                  end
               end
               1081: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[12] ");
                  end
               end
               1082: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[13] ");
                  end
               end
               1083: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[14] ");
                  end
               end
               1084: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[15] ");
                  end
               end
               1085: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[16] ");
                  end
               end
               1086: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[17] ");
                  end
               end
               1087: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[18] ");
                  end
               end
               1088: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[19] ");
                  end
               end
               1089: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[20] ");
                  end
               end
               1090: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[21] ");
                  end
               end
               1091: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[22] ");
                  end
               end
               1092: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[23] ");
                  end
               end
               1093: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[24] ");
                  end
               end
               1094: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.COUNTER_CTRL_reg.DR[25] ");
                  end
               end
               1095: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.SIB_CBB.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1096: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.CBB_reg.DR[27:0], load value = 1111000000001111111111111111");
               end
               1097: begin
                  $display($realtime, "ns:   u_upm_2.upm_inst.CBB_reg.DR[27:0], expected value = 1111000000001111111111111111");
               end
               1098: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[0] ");
                  end
               end
               1099: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[1] ");
                  end
               end
               1100: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[2] ");
                  end
               end
               1101: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[3] ");
                  end
               end
               1102: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[4] ");
                  end
               end
               1103: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[5] ");
                  end
               end
               1104: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[6] ");
                  end
               end
               1105: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[7] ");
                  end
               end
               1106: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[8] ");
                  end
               end
               1107: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[9] ");
                  end
               end
               1108: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[10] ");
                  end
               end
               1109: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[11] ");
                  end
               end
               1110: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[12] ");
                  end
               end
               1111: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[13] ");
                  end
               end
               1112: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[14] ");
                  end
               end
               1113: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[15] ");
                  end
               end
               1114: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[16] ");
                  end
               end
               1115: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[17] ");
                  end
               end
               1116: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[18] ");
                  end
               end
               1117: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[19] ");
                  end
               end
               1118: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[20] ");
                  end
               end
               1119: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[21] ");
                  end
               end
               1120: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[22] ");
                  end
               end
               1121: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[23] ");
                  end
               end
               1122: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[24] ");
                  end
               end
               1123: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[25] ");
                  end
               end
               1124: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[26] ");
                  end
               end
               1125: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_2.upm_inst.CBB_reg.DR[27] ");
                  end
               end
               1126: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_UPM_STATUS.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1127: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.UPM_STATUS_reg.DR[24:0], load value = 1110000000011111111111111");
               end
               1128: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.UPM_STATUS_reg.DR[24:0], expected value = 1110000000011111111111111");
               end
               1129: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[0] ");
                  end
               end
               1130: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[1] ");
                  end
               end
               1131: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[2] ");
                  end
               end
               1132: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[3] ");
                  end
               end
               1133: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[4] ");
                  end
               end
               1134: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[5] ");
                  end
               end
               1135: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[6] ");
                  end
               end
               1136: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[7] ");
                  end
               end
               1137: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[8] ");
                  end
               end
               1138: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[9] ");
                  end
               end
               1139: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[10] ");
                  end
               end
               1140: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[11] ");
                  end
               end
               1141: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[12] ");
                  end
               end
               1142: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[13] ");
                  end
               end
               1143: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[14] ");
                  end
               end
               1144: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[15] ");
                  end
               end
               1145: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[16] ");
                  end
               end
               1146: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[17] ");
                  end
               end
               1147: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[18] ");
                  end
               end
               1148: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[19] ");
                  end
               end
               1149: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[20] ");
                  end
               end
               1150: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[21] ");
                  end
               end
               1151: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[22] ");
                  end
               end
               1152: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[23] ");
                  end
               end
               1153: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.UPM_STATUS_reg.DR[24] ");
                  end
               end
               1154: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_RESULT.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1155: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[20:0], load value = 110000000011111111111");
               end
               1156: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[20:0], expected value = 110000000011111111111");
               end
               1157: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[0] ");
                  end
               end
               1158: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[1] ");
                  end
               end
               1159: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[2] ");
                  end
               end
               1160: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[3] ");
                  end
               end
               1161: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[4] ");
                  end
               end
               1162: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[5] ");
                  end
               end
               1163: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[6] ");
                  end
               end
               1164: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[7] ");
                  end
               end
               1165: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[8] ");
                  end
               end
               1166: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[9] ");
                  end
               end
               1167: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[10] ");
                  end
               end
               1168: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[11] ");
                  end
               end
               1169: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[12] ");
                  end
               end
               1170: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[13] ");
                  end
               end
               1171: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[14] ");
                  end
               end
               1172: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[15] ");
                  end
               end
               1173: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[16] ");
                  end
               end
               1174: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[17] ");
                  end
               end
               1175: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[18] ");
                  end
               end
               1176: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[19] ");
                  end
               end
               1177: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_RESULT_reg.DR[20] ");
                  end
               end
               1178: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_COUNTER_CTRL.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1179: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[25:0], load value = 10000000011111111111111110");
               end
               1180: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[25:0], expected value = 10000000011111111111111110");
               end
               1181: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[0] ");
                  end
               end
               1182: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[1] ");
                  end
               end
               1183: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[2] ");
                  end
               end
               1184: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[3] ");
                  end
               end
               1185: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[4] ");
                  end
               end
               1186: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[5] ");
                  end
               end
               1187: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[6] ");
                  end
               end
               1188: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[7] ");
                  end
               end
               1189: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[8] ");
                  end
               end
               1190: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[9] ");
                  end
               end
               1191: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[10] ");
                  end
               end
               1192: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[11] ");
                  end
               end
               1193: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[12] ");
                  end
               end
               1194: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[13] ");
                  end
               end
               1195: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[14] ");
                  end
               end
               1196: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[15] ");
                  end
               end
               1197: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[16] ");
                  end
               end
               1198: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[17] ");
                  end
               end
               1199: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[18] ");
                  end
               end
               1200: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[19] ");
                  end
               end
               1201: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[20] ");
                  end
               end
               1202: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[21] ");
                  end
               end
               1203: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[22] ");
                  end
               end
               1204: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[23] ");
                  end
               end
               1205: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[24] ");
                  end
               end
               1206: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.COUNTER_CTRL_reg.DR[25] ");
                  end
               end
               1207: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.SIB_CBB.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = inst_so");
               end
               1208: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.CBB_reg.DR[27:0], load value = 0000000011111111111111110000");
               end
               1209: begin
                  $display($realtime, "ns:   u_upm_3.upm_inst.CBB_reg.DR[27:0], expected value = 0000000011111111111111110000");
               end
               1210: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[0] ");
                  end
               end
               1211: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[1] ");
                  end
               end
               1212: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[2] ");
                  end
               end
               1213: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[3] ");
                  end
               end
               1214: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[4] ");
                  end
               end
               1215: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[5] ");
                  end
               end
               1216: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[6] ");
                  end
               end
               1217: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[7] ");
                  end
               end
               1218: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[8] ");
                  end
               end
               1219: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[9] ");
                  end
               end
               1220: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[10] ");
                  end
               end
               1221: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[11] ");
                  end
               end
               1222: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[12] ");
                  end
               end
               1223: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[13] ");
                  end
               end
               1224: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[14] ");
                  end
               end
               1225: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[15] ");
                  end
               end
               1226: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[16] ");
                  end
               end
               1227: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[17] ");
                  end
               end
               1228: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[18] ");
                  end
               end
               1229: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[19] ");
                  end
               end
               1230: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[20] ");
                  end
               end
               1231: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[21] ");
                  end
               end
               1232: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[22] ");
                  end
               end
               1233: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[23] ");
                  end
               end
               1234: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[24] ");
                  end
               end
               1235: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[25] ");
                  end
               end
               1236: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[26] ");
                  end
               end
               1237: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = u_upm_3.upm_inst.CBB_reg.DR[27] ");
                  end
               end
               1238: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_pwrmgmt_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               1239: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_array_pwrmgmt_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               1240: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_array_pwrmgmt_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               1241: begin
                  $display($realtime, "ns:   ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[3:0], load value = 1110");
               end
               1242: begin
                  $display($realtime, "ns:   ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[3:0], expected value = 1110");
               end
               1243: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[0] ");
                  end
               end
               1244: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[1] ");
                  end
               end
               1245: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[2] ");
                  end
               end
               1246: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_pwrmgmt_ctrl_hdspsr_inst.tdr[3] ");
                  end
               end
               1247: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_sib_array_trim_fuse_override_inst.scan_in_mux, selection 1: sib = 1'b1 -> scan_in_mux = ijtag_from_so");
               end
               1248: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_array_trim_fuse_override_secure_mux_inst.M1, selection 0: mux_select = 1'b0 -> M1 = mux_in0");
               end
               1249: begin
                  $display($realtime, "ns:   firebird7_in_gate1_tessent_scanmux_array_trim_fuse_override_secure_mux_inst.M1, selection 1: mux_select = 1'b1 -> M1 = mux_in1");
               end
               1250: begin
                  $display($realtime, "ns:   ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[19:0], load value = 11000011111111000000");
               end
               1251: begin
                  $display($realtime, "ns:   ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[19:0], expected value = 11000011111111000000");
               end
               1252: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[0] ");
                  end
               end
               1253: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[1] ");
                  end
               end
               1254: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[2] ");
                  end
               end
               1255: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[3] ");
                  end
               end
               1256: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[4] ");
                  end
               end
               1257: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[5] ");
                  end
               end
               1258: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[6] ");
                  end
               end
               1259: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[7] ");
                  end
               end
               1260: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[8] ");
                  end
               end
               1261: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[9] ");
                  end
               end
               1262: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[10] ");
                  end
               end
               1263: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[11] ");
                  end
               end
               1264: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[12] ");
                  end
               end
               1265: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[13] ");
                  end
               end
               1266: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[14] ");
                  end
               end
               1267: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[15] ");
                  end
               end
               1268: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[16] ");
                  end
               end
               1269: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[17] ");
                  end
               end
               1270: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[18] ");
                  end
               end
               1271: begin
                  if (_found_fail_per_cycle == 1) begin
                    $display($realtime, "ns: Previous scan out : pin ijtag_so , ICL register = ph0_i_firebird7_in_gate1_tessent_tdr_array_trim_fuse_override_ctrl_hdspsr_inst.tdr[19] ");
                  end
               end
               default: begin
                  $display("ERROR: corrupt message index\n");
                  if (_allow_bad_message_index != 1) begin
                     ->before_finish;
                     #0;
                     $finish;
                  end
               end
            endcase // _message_index
         end
         default: begin
            $display("ERROR: corrupt vector number\n");
            ->before_finish;
            #0;
            $finish;
         end
      endcase
   end // if in_range
      else begin
      case (_pat_type)  // _pat_type = vect[6:4]; 
         3'b011:  begin // status message vector
            _message_index = vect[38:7]; 
            case (_message_index)
               0: begin
                  _chain_test_ = 1;
                  _diag_chain_header = 0;
               end
               1: begin
                  if (_pat_num > -1) begin
                    $display("Skipped chain pattern %d\n",_pat_num);
                  end
                  _chain_test_ = 0;
                  _pat_num = -1;
                  $display("End chain test\n");
               end
               3: begin 
                  _end_vec_file_ok = 1;
                  if (_pat_num > -1) begin
                    if (!_chain_test_) begin
                      $display("Skipped pattern %d\n",_pat_num);
                    end
                  end
               end
               4: begin // start of atpg pattern
                  if (_pat_num > -1) begin
                    if (!_chain_test_) begin
                      _skipped_patterns = _skipped_patterns + 1;
                    end
                  end
                  if (_pat_num > -1) begin
                    if (_chain_test_) begin
                      $display("Skipped chain pattern %d\n",_pat_num);
                    end
                    else begin
                      $display("Skipped pattern %d\n",_pat_num);
                    end
                  end
                  _pat_num = _pat_num + 1;
                  _run_testsetup  = 0;
                  _in_testsetup  = 0;
                  if (_end_after_setup  > 0) begin
                    //simulation complete, exit
                    _index = _max_index + 1;
                    _end_vec_file_ok = 1;
                    _end_simulation = 1;
                    _in_range = 0;
                  end
               end
               default: begin
                  // Skip
               end
            endcase // _message_index
         end
         default: begin
            // Skip
         end
      endcase
      end // else !_in_range
   end // index loop
end // file_cnt loop

if (_save_state == 1) begin
  #1;
  mgcdft_save_signal = 1'b1;
//  $display("Writing checkpoint ICLNetwork.v.dat");
//  $save("ICLNetwork.v.dat");
  if (_in_restart == 2) begin
    _in_restart = 1;
  end
  _end_vec_file_ok = do_finish_summary(_end_vec_file_ok);
  #1;
  $stop;
end
end
end  // while _in_restart
 if (_DIAG_file_header == 1) begin
    if (_diag_scan_header==1) begin
      $fwrite(_diag_file, "last_pattern_applied %d\n", _pattern_count);
    end
    $fwrite(_diag_file, "// failing_patterns=%d simulated_patterns=%d", _fail_pattern_cnt, (_pattern_count+1));
    $fwrite(_diag_file, " simulation_time=", $realtime, ";\n");
    $fwrite(_diag_file, "failure_file_end\n");
    $fclose(_diag_file);
 end


#1;
if (_end_vec_file_ok == 0) begin
  $display("ERROR: Pattern file corrupted, simulation aborted\n");
end
_end_vec_file_ok = do_finish_summary(_end_vec_file_ok);
#1;
->before_finish;
#0;
$finish;
end
endmodule
