//------------------------------------------------------------------------------
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2020 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//  Collateral Description:
//  dteg-upm
//
//  Source organization:
//  DTEG Engineering Group (DTEG)
//
//  Support Information:
//  HSD: https://hsdes.intel.com/appstore/article/#/dft_services.bugeco/create
//
//  Revision:
//  DTEG_UPM_2023WW17_FV_1P1_18A
//
//  Module upm_fabric :  < put your functional description here in plain text >
//
//------------------------------------------------------------------------------
///====================================================================================================================
///
/// upm_fabric.sv
///
/// Unit Owner        : dft_build.pl
///
/// Original Author   : Auto-generated by dft_build
///
/// Copyright (c) 2012 Intel Corporation
/// Intel Proprietary
///
///====================================================================================================================
`ifndef UPM_MODULE_UPM_SYSTEM_CBB_PWREN_DECODER
`define UPM_MODULE_UPM_SYSTEM_CBB_PWREN_DECODER
module upm_system_cbb_pwren_decoder 
(
        input   logic [3:0]      system_cbb_pwr_en_in,
        output  logic [15:0]     system_cbb_pwr_en_out
   );
//------------------------------------------------------------------------------------------------------
assign system_cbb_pwr_en_out = 	(system_cbb_pwr_en_in == 4'h0) ?  16'h0000 : 
								(system_cbb_pwr_en_in == 4'h1)	?  16'h0001 :
								(system_cbb_pwr_en_in == 4'h2) ?  16'h0002 :
								(system_cbb_pwr_en_in == 4'h3) ?  16'h0004 :
								(system_cbb_pwr_en_in == 4'h4) ?  16'h0008 :
								(system_cbb_pwr_en_in == 4'h5) ?  16'h0010 :
								(system_cbb_pwr_en_in == 4'h6) ?  16'h0020 :
								(system_cbb_pwr_en_in == 4'h7) ?  16'h0040 :
								(system_cbb_pwr_en_in == 4'h8) ?  16'h0080 :
								(system_cbb_pwr_en_in == 4'h9) ?  16'h0100 :
								(system_cbb_pwr_en_in == 4'hA) ?  16'h0200 :
								(system_cbb_pwr_en_in == 4'hB) ?  16'h0400 :
								(system_cbb_pwr_en_in == 4'hC) ?  16'h0800 :
								(system_cbb_pwr_en_in == 4'hD) ?  16'h1000 :
								(system_cbb_pwr_en_in == 4'hE) ?  16'h2000 :
								(system_cbb_pwr_en_in == 4'hF) ?  16'h4000 : 'b0;
endmodule
`endif
